module mycpu (
  input  wire          aclk,
  input  wire          aresetn,
  input  wire [7:0]    intrpt,
  output wire [3:0]    arid,
  output wire [31:0]   araddr,
  output wire [7:0]    arlen,
  output wire [2:0]    arsize,
  output wire [1:0]    arburst,
  output wire [1:0]    arlock,
  output wire [3:0]    arcache,
  output wire [2:0]    arprot,
  output wire          arvalid,
  input  wire          arready,
  input  wire [3:0]    rid,
  input  wire [31:0]   rdata,
  input  wire [1:0]    rresp,
  input  wire          rlast,
  input  wire          rvalid,
  output wire          rready,
  output wire [3:0]    awid,
  output wire [31:0]   awaddr,
  output wire [7:0]    awlen,
  output wire [2:0]    awsize,
  output wire [1:0]    awburst,
  output wire [1:0]    awlock,
  output wire [3:0]    awcache,
  output wire [2:0]    awprot,
  output wire          awvalid,
  input  wire          awready,
  output wire [3:0]    wid,
  output wire [31:0]   wdata,
  output wire [3:0]    wstrb,
  output wire          wlast,
  output wire          wvalid,
  input  wire          wready,
  input  wire [3:0]    bid,
  input  wire [1:0]    bresp,
  input  wire          bvalid,
  output wire          bready,
  output wire [31:0]   debug0_wb_pc,
  output wire [3:0]    debug0_wb_rf_wen,
  output wire [4:0]    debug0_wb_rf_wnum,
  output wire [31:0]   debug0_wb_rf_wdata,
  output wire [31:0]   DaRAT_val_0,
  output wire [31:0]   DaRAT_val_1,
  output wire [31:0]   DaRAT_val_2,
  output wire [31:0]   DaRAT_val_3,
  output wire [31:0]   DaRAT_val_4,
  output wire [31:0]   DaRAT_val_5,
  output wire [31:0]   DaRAT_val_6,
  output wire [31:0]   DaRAT_val_7,
  output wire [31:0]   DaRAT_val_8,
  output wire [31:0]   DaRAT_val_9,
  output wire [31:0]   DaRAT_val_10,
  output wire [31:0]   DaRAT_val_11,
  output wire [31:0]   DaRAT_val_12,
  output wire [31:0]   DaRAT_val_13,
  output wire [31:0]   DaRAT_val_14,
  output wire [31:0]   DaRAT_val_15,
  output wire [31:0]   DaRAT_val_16,
  output wire [31:0]   DaRAT_val_17,
  output wire [31:0]   DaRAT_val_18,
  output wire [31:0]   DaRAT_val_19,
  output wire [31:0]   DaRAT_val_20,
  output wire [31:0]   DaRAT_val_21,
  output wire [31:0]   DaRAT_val_22,
  output wire [31:0]   DaRAT_val_23,
  output wire [31:0]   DaRAT_val_24,
  output wire [31:0]   DaRAT_val_25,
  output wire [31:0]   DaRAT_val_26,
  output wire [31:0]   DaRAT_val_27,
  output wire [31:0]   DaRAT_val_28,
  output wire [31:0]   DaRAT_val_29,
  output wire [31:0]   DaRAT_val_30,
  output wire [31:0]   DaRAT_val_31,
  input  wire          break_point,
  input  wire          infor_flag,
  input  wire [4:0]    reg_num,
  output wire          ws_valid,
  output wire [31:0]   rf_rdata,
  output wire [7:0]    DifftestBundle_DifftestInstrCommitIndex_0,
  output wire [7:0]    DifftestBundle_DifftestInstrCommitIndex_1,
  output wire [7:0]    DifftestBundle_DifftestInstrCommitIndex_2,
  output wire [7:0]    DifftestBundle_DifftestInstrCommitIndex_3,
  output wire [7:0]    DifftestBundle_DifftestInstrCommitIndex_4,
  output wire          DifftestBundle_DifftestInstrCommitValid_0,
  output wire          DifftestBundle_DifftestInstrCommitValid_1,
  output wire          DifftestBundle_DifftestInstrCommitValid_2,
  output wire          DifftestBundle_DifftestInstrCommitValid_3,
  output wire          DifftestBundle_DifftestInstrCommitValid_4,
  output wire [63:0]   DifftestBundle_DifftestInstrCommitPC_0,
  output wire [63:0]   DifftestBundle_DifftestInstrCommitPC_1,
  output wire [63:0]   DifftestBundle_DifftestInstrCommitPC_2,
  output wire [63:0]   DifftestBundle_DifftestInstrCommitPC_3,
  output wire [63:0]   DifftestBundle_DifftestInstrCommitPC_4,
  output wire [31:0]   DifftestBundle_DifftestInstrCommitInstr_0,
  output wire [31:0]   DifftestBundle_DifftestInstrCommitInstr_1,
  output wire [31:0]   DifftestBundle_DifftestInstrCommitInstr_2,
  output wire [31:0]   DifftestBundle_DifftestInstrCommitInstr_3,
  output wire [31:0]   DifftestBundle_DifftestInstrCommitInstr_4,
  output wire          DifftestBundle_DifftestSkip_0,
  output wire          DifftestBundle_DifftestSkip_1,
  output wire          DifftestBundle_DifftestSkip_2,
  output wire          DifftestBundle_DifftestSkip_3,
  output wire          DifftestBundle_DifftestSkip_4,
  output wire          DifftestBundle_DifftestIsTlbFill_0,
  output wire          DifftestBundle_DifftestIsTlbFill_1,
  output wire          DifftestBundle_DifftestIsTlbFill_2,
  output wire          DifftestBundle_DifftestIsTlbFill_3,
  output wire          DifftestBundle_DifftestIsTlbFill_4,
  output wire [4:0]    DifftestBundle_DifftestTlbFillIndex_0,
  output wire [4:0]    DifftestBundle_DifftestTlbFillIndex_1,
  output wire [4:0]    DifftestBundle_DifftestTlbFillIndex_2,
  output wire [4:0]    DifftestBundle_DifftestTlbFillIndex_3,
  output wire [4:0]    DifftestBundle_DifftestTlbFillIndex_4,
  output wire          DifftestBundle_DifftestIsCount_0,
  output wire          DifftestBundle_DifftestIsCount_1,
  output wire          DifftestBundle_DifftestIsCount_2,
  output wire          DifftestBundle_DifftestIsCount_3,
  output wire          DifftestBundle_DifftestIsCount_4,
  output wire [63:0]   DifftestBundle_DifftestCount_0,
  output wire [63:0]   DifftestBundle_DifftestCount_1,
  output wire [63:0]   DifftestBundle_DifftestCount_2,
  output wire [63:0]   DifftestBundle_DifftestCount_3,
  output wire [63:0]   DifftestBundle_DifftestCount_4,
  output wire          DifftestBundle_DifftestWen_0,
  output wire          DifftestBundle_DifftestWen_1,
  output wire          DifftestBundle_DifftestWen_2,
  output wire          DifftestBundle_DifftestWen_3,
  output wire          DifftestBundle_DifftestWen_4,
  output wire [7:0]    DifftestBundle_DifftestWdest_0,
  output wire [7:0]    DifftestBundle_DifftestWdest_1,
  output wire [7:0]    DifftestBundle_DifftestWdest_2,
  output wire [7:0]    DifftestBundle_DifftestWdest_3,
  output wire [7:0]    DifftestBundle_DifftestWdest_4,
  output wire [63:0]   DifftestBundle_DifftestWdata_0,
  output wire [63:0]   DifftestBundle_DifftestWdata_1,
  output wire [63:0]   DifftestBundle_DifftestWdata_2,
  output wire [63:0]   DifftestBundle_DifftestWdata_3,
  output wire [63:0]   DifftestBundle_DifftestWdata_4,
  output wire          DifftestBundle_DifftestCsrRstat_0,
  output wire          DifftestBundle_DifftestCsrRstat_1,
  output wire          DifftestBundle_DifftestCsrRstat_2,
  output wire          DifftestBundle_DifftestCsrRstat_3,
  output wire          DifftestBundle_DifftestCsrRstat_4,
  output wire [31:0]   DifftestBundle_DifftestCsrData_0,
  output wire [31:0]   DifftestBundle_DifftestCsrData_1,
  output wire [31:0]   DifftestBundle_DifftestCsrData_2,
  output wire [31:0]   DifftestBundle_DifftestCsrData_3,
  output wire [31:0]   DifftestBundle_DifftestCsrData_4,
  output wire          DifftestBundle_DifftestExcpEventExcpValid,
  output wire          DifftestBundle_DifftestExcpEventEret,
  output wire [31:0]   DifftestBundle_DifftestExcpEventIntrNO,
  output wire [31:0]   DifftestBundle_DifftestExcpEventCause,
  output wire [63:0]   DifftestBundle_DifftestExcpEventEPC,
  output wire [31:0]   DifftestBundle_DifftestExcpEventInst,
  output wire          DifftestBundle_DifftestTrapEventValid,
  output wire [7:0]    DifftestBundle_DifftestStoreEventValid,
  output wire [63:0]   DifftestBundle_DifftestStoreEventPAddr,
  output wire [63:0]   DifftestBundle_DifftestStoreEventVAddr,
  output wire [63:0]   DifftestBundle_DifftestStoreEventData,
  output wire [7:0]    DifftestBundle_DifftestLoadEventValid,
  output wire [63:0]   DifftestBundle_DifftestLoadEventPAddr,
  output wire [63:0]   DifftestBundle_DifftestLoadEventVAddr,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateCRMD,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStatePRMD,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateECFG,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateESTAT,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateERA,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateBADV,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateEENTRY,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateTLBIDX,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateTLBEHI,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateTLBELO0,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateTLBELO1,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateASID,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStatePGDL,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStatePGDH,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateSAVE0,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateSAVE1,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateSAVE2,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateSAVE3,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateTID,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateTCFG,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateTVAL,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateTICLR,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateLLBCTL,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateTLBRENTRY,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateDMW0,
  output wire [63:0]   DifftestBundle_DifftestCSRRegStateDMW1,
  output wire [7:0]    DifftestDelayBundle_DifftestInstrCommitIndex_0,
  output wire [7:0]    DifftestDelayBundle_DifftestInstrCommitIndex_1,
  output wire [7:0]    DifftestDelayBundle_DifftestInstrCommitIndex_2,
  output wire [7:0]    DifftestDelayBundle_DifftestInstrCommitIndex_3,
  output wire [7:0]    DifftestDelayBundle_DifftestInstrCommitIndex_4,
  output wire          DifftestDelayBundle_DifftestInstrCommitValid_0,
  output wire          DifftestDelayBundle_DifftestInstrCommitValid_1,
  output wire          DifftestDelayBundle_DifftestInstrCommitValid_2,
  output wire          DifftestDelayBundle_DifftestInstrCommitValid_3,
  output wire          DifftestDelayBundle_DifftestInstrCommitValid_4,
  output wire [63:0]   DifftestDelayBundle_DifftestInstrCommitPC_0,
  output wire [63:0]   DifftestDelayBundle_DifftestInstrCommitPC_1,
  output wire [63:0]   DifftestDelayBundle_DifftestInstrCommitPC_2,
  output wire [63:0]   DifftestDelayBundle_DifftestInstrCommitPC_3,
  output wire [63:0]   DifftestDelayBundle_DifftestInstrCommitPC_4,
  output wire [31:0]   DifftestDelayBundle_DifftestInstrCommitInstr_0,
  output wire [31:0]   DifftestDelayBundle_DifftestInstrCommitInstr_1,
  output wire [31:0]   DifftestDelayBundle_DifftestInstrCommitInstr_2,
  output wire [31:0]   DifftestDelayBundle_DifftestInstrCommitInstr_3,
  output wire [31:0]   DifftestDelayBundle_DifftestInstrCommitInstr_4,
  output wire          DifftestDelayBundle_DifftestSkip_0,
  output wire          DifftestDelayBundle_DifftestSkip_1,
  output wire          DifftestDelayBundle_DifftestSkip_2,
  output wire          DifftestDelayBundle_DifftestSkip_3,
  output wire          DifftestDelayBundle_DifftestSkip_4,
  output wire          DifftestDelayBundle_DifftestIsTlbFill_0,
  output wire          DifftestDelayBundle_DifftestIsTlbFill_1,
  output wire          DifftestDelayBundle_DifftestIsTlbFill_2,
  output wire          DifftestDelayBundle_DifftestIsTlbFill_3,
  output wire          DifftestDelayBundle_DifftestIsTlbFill_4,
  output wire [4:0]    DifftestDelayBundle_DifftestTlbFillIndex_0,
  output wire [4:0]    DifftestDelayBundle_DifftestTlbFillIndex_1,
  output wire [4:0]    DifftestDelayBundle_DifftestTlbFillIndex_2,
  output wire [4:0]    DifftestDelayBundle_DifftestTlbFillIndex_3,
  output wire [4:0]    DifftestDelayBundle_DifftestTlbFillIndex_4,
  output wire          DifftestDelayBundle_DifftestIsCount_0,
  output wire          DifftestDelayBundle_DifftestIsCount_1,
  output wire          DifftestDelayBundle_DifftestIsCount_2,
  output wire          DifftestDelayBundle_DifftestIsCount_3,
  output wire          DifftestDelayBundle_DifftestIsCount_4,
  output wire [63:0]   DifftestDelayBundle_DifftestCount_0,
  output wire [63:0]   DifftestDelayBundle_DifftestCount_1,
  output wire [63:0]   DifftestDelayBundle_DifftestCount_2,
  output wire [63:0]   DifftestDelayBundle_DifftestCount_3,
  output wire [63:0]   DifftestDelayBundle_DifftestCount_4,
  output wire          DifftestDelayBundle_DifftestWen_0,
  output wire          DifftestDelayBundle_DifftestWen_1,
  output wire          DifftestDelayBundle_DifftestWen_2,
  output wire          DifftestDelayBundle_DifftestWen_3,
  output wire          DifftestDelayBundle_DifftestWen_4,
  output wire [7:0]    DifftestDelayBundle_DifftestWdest_0,
  output wire [7:0]    DifftestDelayBundle_DifftestWdest_1,
  output wire [7:0]    DifftestDelayBundle_DifftestWdest_2,
  output wire [7:0]    DifftestDelayBundle_DifftestWdest_3,
  output wire [7:0]    DifftestDelayBundle_DifftestWdest_4,
  output wire [63:0]   DifftestDelayBundle_DifftestWdata_0,
  output wire [63:0]   DifftestDelayBundle_DifftestWdata_1,
  output wire [63:0]   DifftestDelayBundle_DifftestWdata_2,
  output wire [63:0]   DifftestDelayBundle_DifftestWdata_3,
  output wire [63:0]   DifftestDelayBundle_DifftestWdata_4,
  output wire          DifftestDelayBundle_DifftestCsrRstat_0,
  output wire          DifftestDelayBundle_DifftestCsrRstat_1,
  output wire          DifftestDelayBundle_DifftestCsrRstat_2,
  output wire          DifftestDelayBundle_DifftestCsrRstat_3,
  output wire          DifftestDelayBundle_DifftestCsrRstat_4,
  output wire [31:0]   DifftestDelayBundle_DifftestCsrData_0,
  output wire [31:0]   DifftestDelayBundle_DifftestCsrData_1,
  output wire [31:0]   DifftestDelayBundle_DifftestCsrData_2,
  output wire [31:0]   DifftestDelayBundle_DifftestCsrData_3,
  output wire [31:0]   DifftestDelayBundle_DifftestCsrData_4,
  output wire          DifftestDelayBundle_DifftestExcpEventExcpValid,
  output wire          DifftestDelayBundle_DifftestExcpEventEret,
  output wire [31:0]   DifftestDelayBundle_DifftestExcpEventIntrNO,
  output wire [31:0]   DifftestDelayBundle_DifftestExcpEventCause,
  output wire [63:0]   DifftestDelayBundle_DifftestExcpEventEPC,
  output wire [31:0]   DifftestDelayBundle_DifftestExcpEventInst,
  output wire [7:0]    DifftestDelayBundle_DifftestStoreEventValid,
  output wire [63:0]   DifftestDelayBundle_DifftestStoreEventPAddr,
  output wire [63:0]   DifftestDelayBundle_DifftestStoreEventVAddr,
  output wire [63:0]   DifftestDelayBundle_DifftestStoreEventData,
  output wire [7:0]    DifftestDelayBundle_DifftestLoadEventValid,
  output wire [63:0]   DifftestDelayBundle_DifftestLoadEventPAddr,
  output wire [63:0]   DifftestDelayBundle_DifftestLoadEventVAddr,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_0,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_2,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_3,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_4,
  output reg           _zz_DifftestDelayBundle_DifftestInstrCommitValid_0,
  output reg           _zz_DifftestDelayBundle_DifftestInstrCommitValid_1,
  output reg           _zz_DifftestDelayBundle_DifftestInstrCommitValid_2,
  output reg           _zz_DifftestDelayBundle_DifftestInstrCommitValid_3,
  output reg           _zz_DifftestDelayBundle_DifftestInstrCommitValid_4,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_0,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_2,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_3,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_4,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_0,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_2,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_3,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_4,
  output reg           _zz_DifftestDelayBundle_DifftestSkip_0,
  output reg           _zz_DifftestDelayBundle_DifftestSkip_1,
  output reg           _zz_DifftestDelayBundle_DifftestSkip_2,
  output reg           _zz_DifftestDelayBundle_DifftestSkip_3,
  output reg           _zz_DifftestDelayBundle_DifftestSkip_4,
  output reg           _zz_DifftestDelayBundle_DifftestIsTlbFill_0,
  output reg           _zz_DifftestDelayBundle_DifftestIsTlbFill_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsTlbFill_2,
  output reg           _zz_DifftestDelayBundle_DifftestIsTlbFill_3,
  output reg           _zz_DifftestDelayBundle_DifftestIsTlbFill_4,
  output reg  [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_0,
  output reg  [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_1,
  output reg  [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_2,
  output reg  [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_3,
  output reg  [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_4,
  output reg           _zz_DifftestDelayBundle_DifftestIsCount_0,
  output reg           _zz_DifftestDelayBundle_DifftestIsCount_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsCount_2,
  output reg           _zz_DifftestDelayBundle_DifftestIsCount_3,
  output reg           _zz_DifftestDelayBundle_DifftestIsCount_4,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestCount_0,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestCount_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestCount_2,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestCount_3,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestCount_4,
  output reg           _zz_DifftestDelayBundle_DifftestWen_0,
  output reg           _zz_DifftestDelayBundle_DifftestWen_1,
  output reg           _zz_DifftestDelayBundle_DifftestWen_2,
  output reg           _zz_DifftestDelayBundle_DifftestWen_3,
  output reg           _zz_DifftestDelayBundle_DifftestWen_4,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestWdest_0,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestWdest_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestWdest_2,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestWdest_3,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestWdest_4,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestWdata_0,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestWdata_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestWdata_2,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestWdata_3,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestWdata_4,
  output reg           _zz_DifftestDelayBundle_DifftestCsrRstat_0,
  output reg           _zz_DifftestDelayBundle_DifftestCsrRstat_1,
  output reg           _zz_DifftestDelayBundle_DifftestCsrRstat_2,
  output reg           _zz_DifftestDelayBundle_DifftestCsrRstat_3,
  output reg           _zz_DifftestDelayBundle_DifftestCsrRstat_4,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_0,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_2,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_3,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_4,
  output reg           _zz_DifftestDelayBundle_DifftestExcpEventExcpValid,
  output reg           _zz_DifftestDelayBundle_DifftestExcpEventEret,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestExcpEventIntrNO,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestExcpEventCause,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestExcpEventEPC,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestExcpEventInst,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestStoreEventValid,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestStoreEventPAddr,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestStoreEventVAddr,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestStoreEventData,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestLoadEventValid,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestLoadEventPAddr,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestLoadEventVAddr,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_0_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_1_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_2_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_3_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_4_1,
  output reg           _zz_DifftestDelayBundle_DifftestInstrCommitValid_0_1,
  output reg           _zz_DifftestDelayBundle_DifftestInstrCommitValid_1_1,
  output reg           _zz_DifftestDelayBundle_DifftestInstrCommitValid_2_1,
  output reg           _zz_DifftestDelayBundle_DifftestInstrCommitValid_3_1,
  output reg           _zz_DifftestDelayBundle_DifftestInstrCommitValid_4_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_0_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_1_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_2_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_3_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_4_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_0_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_1_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_2_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_3_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_4_1,
  output reg           _zz_DifftestDelayBundle_DifftestSkip_0_1,
  output reg           _zz_DifftestDelayBundle_DifftestSkip_1_1,
  output reg           _zz_DifftestDelayBundle_DifftestSkip_2_1,
  output reg           _zz_DifftestDelayBundle_DifftestSkip_3_1,
  output reg           _zz_DifftestDelayBundle_DifftestSkip_4_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsTlbFill_0_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsTlbFill_1_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsTlbFill_2_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsTlbFill_3_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsTlbFill_4_1,
  output reg  [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_0_1,
  output reg  [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_1_1,
  output reg  [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_2_1,
  output reg  [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_3_1,
  output reg  [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_4_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsCount_0_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsCount_1_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsCount_2_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsCount_3_1,
  output reg           _zz_DifftestDelayBundle_DifftestIsCount_4_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestCount_0_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestCount_1_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestCount_2_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestCount_3_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestCount_4_1,
  output reg           _zz_DifftestDelayBundle_DifftestWen_0_1,
  output reg           _zz_DifftestDelayBundle_DifftestWen_1_1,
  output reg           _zz_DifftestDelayBundle_DifftestWen_2_1,
  output reg           _zz_DifftestDelayBundle_DifftestWen_3_1,
  output reg           _zz_DifftestDelayBundle_DifftestWen_4_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestWdest_0_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestWdest_1_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestWdest_2_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestWdest_3_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestWdest_4_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestWdata_0_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestWdata_1_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestWdata_2_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestWdata_3_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestWdata_4_1,
  output reg           _zz_DifftestDelayBundle_DifftestCsrRstat_0_1,
  output reg           _zz_DifftestDelayBundle_DifftestCsrRstat_1_1,
  output reg           _zz_DifftestDelayBundle_DifftestCsrRstat_2_1,
  output reg           _zz_DifftestDelayBundle_DifftestCsrRstat_3_1,
  output reg           _zz_DifftestDelayBundle_DifftestCsrRstat_4_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_0_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_1_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_2_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_3_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_4_1,
  output reg           _zz_DifftestDelayBundle_DifftestExcpEventExcpValid_1,
  output reg           _zz_DifftestDelayBundle_DifftestExcpEventEret_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestExcpEventIntrNO_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestExcpEventCause_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestExcpEventEPC_1,
  output reg  [31:0]   _zz_DifftestDelayBundle_DifftestExcpEventInst_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestStoreEventValid_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestStoreEventPAddr_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestStoreEventVAddr_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestStoreEventData_1,
  output reg  [7:0]    _zz_DifftestDelayBundle_DifftestLoadEventValid_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestLoadEventPAddr_1,
  output reg  [63:0]   _zz_DifftestDelayBundle_DifftestLoadEventVAddr_1
);
  localparam ALUOp_add = 4'd0;
  localparam ALUOp_sub = 4'd1;
  localparam ALUOp_slt = 4'd2;
  localparam ALUOp_sltu = 4'd3;
  localparam ALUOp_eq = 4'd4;
  localparam ALUOp_nor_1 = 4'd5;
  localparam ALUOp_and_1 = 4'd6;
  localparam ALUOp_or_1 = 4'd7;
  localparam ALUOp_xor_1 = 4'd8;
  localparam ALUOp_sll_1 = 4'd9;
  localparam ALUOp_srl_1 = 4'd10;
  localparam ALUOp_sra_1 = 4'd11;
  localparam ALUOp_passa = 4'd12;
  localparam ALUOp_passb = 4'd13;
  localparam BRUOp_nop = 2'd0;
  localparam BRUOp_add = 2'd1;
  localparam BRUOp_cadd = 2'd2;
  localparam BRUOp_ncadd = 2'd3;
  localparam CRUOp_nop = 2'd0;
  localparam CRUOp_pass = 2'd1;
  localparam CRUOp_mask = 2'd2;
  localparam ALUROOp_reg_1 = 3'd0;
  localparam ALUROOp_regimm = 3'd1;
  localparam ALUROOp_pcimm = 3'd2;
  localparam ALUROOp_csr = 3'd3;
  localparam ALUROOp_linkpc = 3'd4;
  localparam ALUROOp_linkreg = 3'd5;
  localparam CRUROOp_id = 2'd0;
  localparam CRUROOp_lo = 2'd1;
  localparam CRUROOp_hi = 2'd2;
  localparam MULUOp_mullo = 2'd0;
  localparam MULUOp_mulhi = 2'd1;
  localparam MULUOp_mulhiu = 2'd2;
  localparam DIVUOp_div = 2'd0;
  localparam DIVUOp_divu = 2'd1;
  localparam DIVUOp_mod_1 = 2'd2;
  localparam DIVUOp_modu = 2'd3;
  localparam LSUOp_cacop = 4'd0;
  localparam LSUOp_tlbsrch = 4'd1;
  localparam LSUOp_tlbrd = 4'd2;
  localparam LSUOp_tlbwr = 4'd3;
  localparam LSUOp_tlbfill = 4'd4;
  localparam LSUOp_invtlb = 4'd5;
  localparam LSUOp_ll = 4'd6;
  localparam LSUOp_sc = 4'd7;
  localparam LSUOp_ld = 4'd8;
  localparam LSUOp_ldu = 4'd9;
  localparam LSUOp_st = 4'd10;
  localparam LSUOp_preld = 4'd11;
  localparam LSUOp_dbar = 4'd12;
  localparam LSUOp_ibar = 4'd13;
  localparam LSUROOp_reg_1 = 1'd0;
  localparam LSUROOp_regimm = 1'd1;
  localparam TLBOp_nop = 3'd0;
  localparam TLBOp_srch = 3'd1;
  localparam TLBOp_read = 3'd2;
  localparam TLBOp_write = 3'd3;
  localparam TLBOp_fill = 3'd4;
  localparam TLBOp_inv = 3'd5;
  localparam ROBSpecialOp_nop = 4'd0;
  localparam ROBSpecialOp_bpuUpdate = 4'd1;
  localparam ROBSpecialOp_lsuAction = 4'd2;
  localparam ROBSpecialOp_ll = 4'd3;
  localparam ROBSpecialOp_writeCSR = 4'd4;
  localparam ROBSpecialOp_ertn = 4'd5;
  localparam ROBSpecialOp_idle = 4'd6;
  localparam ROBSpecialOp_readCSR = 4'd7;
  localparam ROBSpecialOp_readCNT = 4'd8;
  localparam LSUSizeOp_byte_1 = 4'd1;
  localparam LSUSizeOp_halfword = 4'd3;
  localparam LSUSizeOp_word = 4'd15;
  localparam FUType_alu = 3'd0;
  localparam FUType_csr = 3'd1;
  localparam FUType_counter = 3'd2;
  localparam FUType_lsu = 3'd3;
  localparam FUType_mulu = 3'd4;
  localparam FUType_divu = 3'd5;

  reg                 cpuClockingArea_fuLSU_io_output_ready;
  reg                 cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_ready;
  reg                 cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_ready;
  reg                 cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_ready;
  reg                 cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_ready;
  reg                 cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_ready;
  reg                 cpuClockingArea_areaFlushReset_roALU0_io_toFU_ready;
  reg                 cpuClockingArea_areaFlushReset_roALU1_io_toFU_ready;
  reg                 cpuClockingArea_areaFlushReset_roMULU_io_toFU_ready;
  reg                 cpuClockingArea_areaFlushReset_roDIVU_io_toFU_ready;
  reg                 cpuClockingArea_areaFlushReset_roLSU_io_toFU_ready;
  reg                 cpuClockingArea_areaFlushReset_fuALU0_io_output_ready;
  reg                 cpuClockingArea_areaFlushReset_fuALU1_io_output_ready;
  reg                 cpuClockingArea_areaFlushReset_fuMULU_io_output_ready;
  reg                 cpuClockingArea_areaFlushReset_fuDIVU_io_output_ready;
  wire       [3:0]    cpuClockingArea_arbiter_io_out_arid;
  wire       [31:0]   cpuClockingArea_arbiter_io_out_araddr;
  wire       [7:0]    cpuClockingArea_arbiter_io_out_arlen;
  wire       [2:0]    cpuClockingArea_arbiter_io_out_arsize;
  wire       [1:0]    cpuClockingArea_arbiter_io_out_arburst;
  wire       [1:0]    cpuClockingArea_arbiter_io_out_arlock;
  wire       [3:0]    cpuClockingArea_arbiter_io_out_arcache;
  wire       [2:0]    cpuClockingArea_arbiter_io_out_arprot;
  wire                cpuClockingArea_arbiter_io_out_arvalid;
  wire                cpuClockingArea_arbiter_io_out_rready;
  wire       [3:0]    cpuClockingArea_arbiter_io_out_awid;
  wire       [31:0]   cpuClockingArea_arbiter_io_out_awaddr;
  wire       [7:0]    cpuClockingArea_arbiter_io_out_awlen;
  wire       [2:0]    cpuClockingArea_arbiter_io_out_awsize;
  wire       [1:0]    cpuClockingArea_arbiter_io_out_awburst;
  wire       [1:0]    cpuClockingArea_arbiter_io_out_awlock;
  wire       [3:0]    cpuClockingArea_arbiter_io_out_awcache;
  wire       [2:0]    cpuClockingArea_arbiter_io_out_awprot;
  wire                cpuClockingArea_arbiter_io_out_awvalid;
  wire       [3:0]    cpuClockingArea_arbiter_io_out_wid;
  wire       [31:0]   cpuClockingArea_arbiter_io_out_wdata;
  wire       [3:0]    cpuClockingArea_arbiter_io_out_wstrb;
  wire                cpuClockingArea_arbiter_io_out_wlast;
  wire                cpuClockingArea_arbiter_io_out_wvalid;
  wire                cpuClockingArea_arbiter_io_out_bready;
  wire                cpuClockingArea_arbiter_io_iCache_arready;
  wire       [3:0]    cpuClockingArea_arbiter_io_iCache_rid;
  wire       [31:0]   cpuClockingArea_arbiter_io_iCache_rdata;
  wire       [1:0]    cpuClockingArea_arbiter_io_iCache_rresp;
  wire                cpuClockingArea_arbiter_io_iCache_rlast;
  wire                cpuClockingArea_arbiter_io_iCache_rvalid;
  wire                cpuClockingArea_arbiter_io_dCache_arready;
  wire       [3:0]    cpuClockingArea_arbiter_io_dCache_rid;
  wire       [31:0]   cpuClockingArea_arbiter_io_dCache_rdata;
  wire       [1:0]    cpuClockingArea_arbiter_io_dCache_rresp;
  wire                cpuClockingArea_arbiter_io_dCache_rlast;
  wire                cpuClockingArea_arbiter_io_dCache_rvalid;
  wire                cpuClockingArea_arbiter_io_dCache_awready;
  wire                cpuClockingArea_arbiter_io_dCache_wready;
  wire       [3:0]    cpuClockingArea_arbiter_io_dCache_bid;
  wire       [1:0]    cpuClockingArea_arbiter_io_dCache_bresp;
  wire                cpuClockingArea_arbiter_io_dCache_bvalid;
  wire                cpuClockingArea_tlb_io_iCacheReq_hit;
  wire       [19:0]   cpuClockingArea_tlb_io_iCacheReq_pageInfo_ppn;
  wire       [1:0]    cpuClockingArea_tlb_io_iCacheReq_pageInfo_plv;
  wire       [1:0]    cpuClockingArea_tlb_io_iCacheReq_pageInfo_mat;
  wire                cpuClockingArea_tlb_io_iCacheReq_pageInfo_d;
  wire                cpuClockingArea_tlb_io_iCacheReq_pageInfo_v;
  wire                cpuClockingArea_tlb_io_dCacheReq_hit;
  wire       [19:0]   cpuClockingArea_tlb_io_dCacheReq_pageInfo_ppn;
  wire       [1:0]    cpuClockingArea_tlb_io_dCacheReq_pageInfo_plv;
  wire       [1:0]    cpuClockingArea_tlb_io_dCacheReq_pageInfo_mat;
  wire                cpuClockingArea_tlb_io_dCacheReq_pageInfo_d;
  wire                cpuClockingArea_tlb_io_dCacheReq_pageInfo_v;
  wire       [1:0]    cpuClockingArea_tlb__zz_io_swRead_value_2;
  wire       [21:0]   cpuClockingArea_tlb__zz_io_swRead_value_3;
  wire       [5:0]    cpuClockingArea_tlb__zz_io_swRead_value_4;
  wire                cpuClockingArea_tlb__zz_io_swRead_value_5;
  wire                cpuClockingArea_tlb__zz_io_swRead_value_6;
  wire       [12:0]   cpuClockingArea_tlb__zz_io_swRead_value_7;
  wire       [18:0]   cpuClockingArea_tlb__zz_io_swRead_value_8;
  wire                cpuClockingArea_tlb__zz_io_swRead_value_9;
  wire                cpuClockingArea_tlb__zz_io_swRead_value_10;
  wire       [1:0]    cpuClockingArea_tlb__zz_io_swRead_value_11;
  wire       [1:0]    cpuClockingArea_tlb__zz_io_swRead_value_12;
  wire                cpuClockingArea_tlb__zz_io_swRead_value_13;
  wire                cpuClockingArea_tlb__zz_io_swRead_value_14;
  wire       [19:0]   cpuClockingArea_tlb__zz_io_swRead_value_15;
  wire       [3:0]    cpuClockingArea_tlb__zz_io_swRead_value_16;
  wire                cpuClockingArea_tlb__zz_io_swRead_value_17;
  wire                cpuClockingArea_tlb__zz_io_swRead_value_18;
  wire       [1:0]    cpuClockingArea_tlb__zz_io_swRead_value_19;
  wire       [1:0]    cpuClockingArea_tlb__zz_io_swRead_value_20;
  wire                cpuClockingArea_tlb__zz_io_swRead_value_21;
  wire                cpuClockingArea_tlb__zz_io_swRead_value_22;
  wire       [19:0]   cpuClockingArea_tlb__zz_io_swRead_value_23;
  wire       [3:0]    cpuClockingArea_tlb__zz_io_swRead_value_24;
  wire       [9:0]    cpuClockingArea_tlb_io_csrWrite_asid;
  wire                cpuClockingArea_tlb_io_csrWrite_idxWen;
  wire                cpuClockingArea_tlb_io_csrWrite_entryWen;
  wire                cpuClockingArea_memService_io_iCacheCtrl_stall;
  wire       [31:0]   cpuClockingArea_memService_io_iCacheCtrl_cacopVA;
  wire                cpuClockingArea_memService_io_iCacheCtrl_cacopStoreTag;
  wire                cpuClockingArea_memService_io_iCacheCtrl_cacopIndexInvalidate;
  wire                cpuClockingArea_memService_io_iCacheCtrl_cacopHitInvalidate;
  wire                cpuClockingArea_memService_io_dCacheCtrl_stall;
  wire       [31:0]   cpuClockingArea_memService_io_dCacheCtrl_cacopVA;
  wire                cpuClockingArea_memService_io_dCacheCtrl_cacopStoreTag;
  wire                cpuClockingArea_memService_io_dCacheCtrl_cacopIndexInvalidate;
  wire                cpuClockingArea_memService_io_dCacheCtrl_cacopHitInvalidate;
  wire       [2:0]    cpuClockingArea_memService_io_TLBCtrl_op;
  wire                cpuClockingArea_memService_io_TLBCtrl_invGlobal;
  wire                cpuClockingArea_memService_io_TLBCtrl_invLocal;
  wire                cpuClockingArea_memService_io_TLBCtrl_invLocalVAMatch;
  wire                cpuClockingArea_memService_io_TLBCtrl_invLocalVANotMatch;
  wire       [1:0]    cpuClockingArea_memService_io_TLBCtrl_index;
  wire       [18:0]   cpuClockingArea_memService_io_TLBCtrl_invVA;
  wire       [9:0]    cpuClockingArea_memService_io_TLBCtrl_asid;
  wire       [5:0]    cpuClockingArea_sRAT_io_srcReadPort_0_0_prd;
  wire                cpuClockingArea_sRAT_io_srcReadPort_0_0_valid;
  wire       [5:0]    cpuClockingArea_sRAT_io_srcReadPort_0_1_prd;
  wire                cpuClockingArea_sRAT_io_srcReadPort_0_1_valid;
  wire       [5:0]    cpuClockingArea_sRAT_io_srcReadPort_1_0_prd;
  wire                cpuClockingArea_sRAT_io_srcReadPort_1_0_valid;
  wire       [5:0]    cpuClockingArea_sRAT_io_srcReadPort_1_1_prd;
  wire                cpuClockingArea_sRAT_io_srcReadPort_1_1_valid;
  wire       [5:0]    cpuClockingArea_sRAT_io_prevPRDReadPort_0_prd;
  wire                cpuClockingArea_sRAT_io_prevPRDReadPort_0_valid;
  wire       [5:0]    cpuClockingArea_sRAT_io_prevPRDReadPort_1_prd;
  wire                cpuClockingArea_sRAT_io_prevPRDReadPort_1_valid;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_0;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_1;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_2;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_3;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_4;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_5;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_6;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_7;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_8;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_9;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_10;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_11;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_12;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_13;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_14;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_15;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_16;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_17;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_18;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_19;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_20;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_21;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_22;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_23;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_24;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_25;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_26;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_27;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_28;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_29;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_30;
  wire       [5:0]    cpuClockingArea_aRAT_io_recoveryPort_31;
  wire       [1:0]    cpuClockingArea_freeList_io_dispatch_availMask;
  wire       [5:0]    cpuClockingArea_freeList_io_dispatch_prfIdx_0;
  wire       [5:0]    cpuClockingArea_freeList_io_dispatch_prfIdx_1;
  wire                cpuClockingArea_pc_io_iCacheFeed_0_valid;
  wire       [31:0]   cpuClockingArea_pc_io_iCacheFeed_0_payload_address;
  wire       [3:0]    cpuClockingArea_pc_io_iCacheFeed_0_payload_size;
  wire       [31:0]   cpuClockingArea_pc_io_iCacheFeed_0_payload_branchInfo_predictPC;
  wire                cpuClockingArea_pc_io_iCacheFeed_0_payload_branchInfo_predictResult;
  wire                cpuClockingArea_pc_io_iCacheFeed_1_valid;
  wire       [31:0]   cpuClockingArea_pc_io_iCacheFeed_1_payload_address;
  wire       [3:0]    cpuClockingArea_pc_io_iCacheFeed_1_payload_size;
  wire       [31:0]   cpuClockingArea_pc_io_iCacheFeed_1_payload_branchInfo_predictPC;
  wire                cpuClockingArea_pc_io_iCacheFeed_1_payload_branchInfo_predictResult;
  wire                cpuClockingArea_pc_io_pc_0_valid;
  wire       [31:0]   cpuClockingArea_pc_io_pc_0_payload;
  wire                cpuClockingArea_pc_io_pc_1_valid;
  wire       [31:0]   cpuClockingArea_pc_io_pc_1_payload;
  wire                cpuClockingArea_nextLinePredictor_io_npc_0_valid;
  wire       [31:0]   cpuClockingArea_nextLinePredictor_io_npc_0_payload;
  wire                cpuClockingArea_nextLinePredictor_io_npc_1_valid;
  wire       [31:0]   cpuClockingArea_nextLinePredictor_io_npc_1_payload;
  wire       [31:0]   cpuClockingArea_nextLinePredictor_io_branchInfo_0_predictPC;
  wire                cpuClockingArea_nextLinePredictor_io_branchInfo_0_predictResult;
  wire       [31:0]   cpuClockingArea_nextLinePredictor_io_branchInfo_1_predictPC;
  wire                cpuClockingArea_nextLinePredictor_io_branchInfo_1_predictResult;
  wire                cpuClockingArea_iCache_io_input_0_ready;
  wire                cpuClockingArea_iCache_io_input_1_ready;
  wire       [1:0]    cpuClockingArea_iCache_io_output_availMask;
  wire       [31:0]   cpuClockingArea_iCache_io_output_info_0_inst;
  wire       [31:0]   cpuClockingArea_iCache_io_output_info_0_branchInfo_predictPC;
  wire                cpuClockingArea_iCache_io_output_info_0_branchInfo_predictResult;
  wire                cpuClockingArea_iCache_io_output_info_0_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_iCache_io_output_info_0_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_iCache_io_output_info_0_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_iCache_io_output_info_0_pc;
  wire       [31:0]   cpuClockingArea_iCache_io_output_info_1_inst;
  wire       [31:0]   cpuClockingArea_iCache_io_output_info_1_branchInfo_predictPC;
  wire                cpuClockingArea_iCache_io_output_info_1_branchInfo_predictResult;
  wire                cpuClockingArea_iCache_io_output_info_1_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_iCache_io_output_info_1_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_iCache_io_output_info_1_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_iCache_io_output_info_1_pc;
  wire       [19:0]   cpuClockingArea_iCache_io_tlb_virtPageNumber;
  wire                cpuClockingArea_iCache_io_ctrl_busy;
  wire       [31:0]   cpuClockingArea_iCache_io_badv_vaddr;
  wire                cpuClockingArea_iCache_io_badv_wen;
  wire       [3:0]    cpuClockingArea_iCache_io_axi_arid;
  wire       [31:0]   cpuClockingArea_iCache_io_axi_araddr;
  wire       [7:0]    cpuClockingArea_iCache_io_axi_arlen;
  wire       [2:0]    cpuClockingArea_iCache_io_axi_arsize;
  wire       [1:0]    cpuClockingArea_iCache_io_axi_arburst;
  wire       [1:0]    cpuClockingArea_iCache_io_axi_arlock;
  wire       [3:0]    cpuClockingArea_iCache_io_axi_arcache;
  wire       [2:0]    cpuClockingArea_iCache_io_axi_arprot;
  wire                cpuClockingArea_iCache_io_axi_arvalid;
  wire                cpuClockingArea_iCache_io_axi_rready;
  wire                cpuClockingArea_fuLSU_io_input_ready;
  wire                cpuClockingArea_fuLSU_io_output_valid;
  wire       [4:0]    cpuClockingArea_fuLSU_io_output_payload_robIdx;
  wire       [31:0]   cpuClockingArea_fuLSU_io_output_payload_data;
  wire       [5:0]    cpuClockingArea_fuLSU_io_output_payload_prd;
  wire       [31:0]   cpuClockingArea_fuLSU_io_output_payload_branchResult_targetPC;
  wire                cpuClockingArea_fuLSU_io_output_payload_branchResult_branchResult;
  wire                cpuClockingArea_fuLSU_io_output_payload_branchResult_predictFail;
  wire                cpuClockingArea_fuLSU_io_output_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_fuLSU_io_output_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_fuLSU_io_output_payload_exceptionInfo_eSubCode;
  wire                cpuClockingArea_fuLSU_io_wakeOut_0_valid;
  wire       [5:0]    cpuClockingArea_fuLSU_io_wakeOut_0_payload;
  wire                cpuClockingArea_fuLSU_io_wakeOut_1_valid;
  wire       [5:0]    cpuClockingArea_fuLSU_io_wakeOut_1_payload;
  wire       [19:0]   cpuClockingArea_fuLSU_io_tlb_virtPageNumber;
  wire       [31:0]   cpuClockingArea_fuLSU_io_llBitComm_toUpdateAddr;
  wire                cpuClockingArea_fuLSU_io_llBitComm_wen;
  wire                cpuClockingArea_fuLSU_io_ctrl_busy;
  wire                cpuClockingArea_fuLSU_io_specialOpBufferUpdate_valid;
  wire       [3:0]    cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_uop_lsuOp;
  wire       [4:0]    cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_uop_lsuCoOp;
  wire       [31:0]   cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_vaddr;
  wire       [9:0]    cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_asid;
  wire       [4:0]    cpuClockingArea_fuLSU_io_badv_robIdx;
  wire       [31:0]   cpuClockingArea_fuLSU_io_badv_vaddr;
  wire                cpuClockingArea_fuLSU_io_badv_wen;
  wire       [3:0]    cpuClockingArea_fuLSU_io_axi_arid;
  wire       [31:0]   cpuClockingArea_fuLSU_io_axi_araddr;
  wire       [7:0]    cpuClockingArea_fuLSU_io_axi_arlen;
  wire       [2:0]    cpuClockingArea_fuLSU_io_axi_arsize;
  wire       [1:0]    cpuClockingArea_fuLSU_io_axi_arburst;
  wire       [1:0]    cpuClockingArea_fuLSU_io_axi_arlock;
  wire       [3:0]    cpuClockingArea_fuLSU_io_axi_arcache;
  wire       [2:0]    cpuClockingArea_fuLSU_io_axi_arprot;
  wire                cpuClockingArea_fuLSU_io_axi_arvalid;
  wire                cpuClockingArea_fuLSU_io_axi_rready;
  wire       [3:0]    cpuClockingArea_fuLSU_io_axi_awid;
  wire       [31:0]   cpuClockingArea_fuLSU_io_axi_awaddr;
  wire       [7:0]    cpuClockingArea_fuLSU_io_axi_awlen;
  wire       [2:0]    cpuClockingArea_fuLSU_io_axi_awsize;
  wire       [1:0]    cpuClockingArea_fuLSU_io_axi_awburst;
  wire       [1:0]    cpuClockingArea_fuLSU_io_axi_awlock;
  wire       [3:0]    cpuClockingArea_fuLSU_io_axi_awcache;
  wire       [2:0]    cpuClockingArea_fuLSU_io_axi_awprot;
  wire                cpuClockingArea_fuLSU_io_axi_awvalid;
  wire       [3:0]    cpuClockingArea_fuLSU_io_axi_wid;
  wire       [31:0]   cpuClockingArea_fuLSU_io_axi_wdata;
  wire       [3:0]    cpuClockingArea_fuLSU_io_axi_wstrb;
  wire                cpuClockingArea_fuLSU_io_axi_wlast;
  wire                cpuClockingArea_fuLSU_io_axi_wvalid;
  wire                cpuClockingArea_fuLSU_io_axi_bready;
  wire       [31:0]   cpuClockingArea_fuLSU_io_storeData;
  wire       [3:0]    cpuClockingArea_fuLSU_io_storeMask;
  wire       [3:0]    cpuClockingArea_fuLSU_io_loadMask;
  wire       [31:0]   cpuClockingArea_fuLSU_io_VAddr;
  wire       [31:0]   cpuClockingArea_fuLSU_io_PAddr;
  wire       [31:0]   cpuClockingArea_prf_io_read_0_0_data;
  wire       [31:0]   cpuClockingArea_prf_io_read_0_1_data;
  wire       [31:0]   cpuClockingArea_prf_io_read_1_0_data;
  wire       [31:0]   cpuClockingArea_prf_io_read_1_1_data;
  wire       [31:0]   cpuClockingArea_prf_io_read_2_0_data;
  wire       [31:0]   cpuClockingArea_prf_io_read_2_1_data;
  wire       [31:0]   cpuClockingArea_prf_io_read_3_0_data;
  wire       [31:0]   cpuClockingArea_prf_io_read_3_1_data;
  wire       [31:0]   cpuClockingArea_prf_io_read_4_0_data;
  wire       [31:0]   cpuClockingArea_prf_io_read_4_1_data;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_0;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_1;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_2;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_3;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_4;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_5;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_6;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_7;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_8;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_9;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_10;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_11;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_12;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_13;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_14;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_15;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_16;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_17;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_18;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_19;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_20;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_21;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_22;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_23;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_24;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_25;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_26;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_27;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_28;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_29;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_30;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_31;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_32;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_33;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_34;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_35;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_36;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_37;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_38;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_39;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_40;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_41;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_42;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_43;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_44;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_45;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_46;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_47;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_48;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_49;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_50;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_51;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_52;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_53;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_54;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_55;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_56;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_57;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_58;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_59;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_60;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_61;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_62;
  wire       [31:0]   cpuClockingArea_prf_io_debugRegs_63;
  wire       [1:0]    cpuClockingArea_rob_io_dispatch_availMask;
  wire       [4:0]    cpuClockingArea_rob_io_dispatch_robIdx_0;
  wire       [4:0]    cpuClockingArea_rob_io_dispatch_robIdx_1;
  wire       [5:0]    cpuClockingArea_rob_io_retireARAT_0_prd;
  wire       [4:0]    cpuClockingArea_rob_io_retireARAT_0_ard;
  wire                cpuClockingArea_rob_io_retireARAT_0_wen;
  wire       [5:0]    cpuClockingArea_rob_io_retireARAT_1_prd;
  wire       [4:0]    cpuClockingArea_rob_io_retireARAT_1_ard;
  wire                cpuClockingArea_rob_io_retireARAT_1_wen;
  wire       [5:0]    cpuClockingArea_rob_io_retireFreeList_prfIdx_0;
  wire       [5:0]    cpuClockingArea_rob_io_retireFreeList_prfIdx_1;
  wire       [1:0]    cpuClockingArea_rob_io_retireFreeList_writeNum;
  wire                cpuClockingArea_rob_io_retireFreeList_delayedFlush;
  wire       [4:0]    cpuClockingArea_rob_io_retireLSU_robIdx_0;
  wire       [4:0]    cpuClockingArea_rob_io_retireLSU_robIdx_1;
  wire                cpuClockingArea_rob_io_retireLSU_allowRetire_0;
  wire                cpuClockingArea_rob_io_retireLSU_allowRetire_1;
  wire                cpuClockingArea_rob_io_wakeupMem;
  wire                cpuClockingArea_rob_io_updateBPU_0_valid;
  wire       [31:0]   cpuClockingArea_rob_io_updateBPU_0_payload_pc;
  wire                cpuClockingArea_rob_io_updateBPU_0_payload_isJumpInst;
  wire                cpuClockingArea_rob_io_updateBPU_0_payload_taken;
  wire                cpuClockingArea_rob_io_updateBPU_0_payload_predictFail;
  wire       [31:0]   cpuClockingArea_rob_io_updateBPU_0_payload_target;
  wire                cpuClockingArea_rob_io_updateBPU_1_valid;
  wire       [31:0]   cpuClockingArea_rob_io_updateBPU_1_payload_pc;
  wire                cpuClockingArea_rob_io_updateBPU_1_payload_isJumpInst;
  wire                cpuClockingArea_rob_io_updateBPU_1_payload_taken;
  wire                cpuClockingArea_rob_io_updateBPU_1_payload_predictFail;
  wire       [31:0]   cpuClockingArea_rob_io_updateBPU_1_payload_target;
  wire                cpuClockingArea_rob_io_csrCtrl_llBitUpdate;
  wire                cpuClockingArea_rob_io_csrCtrl_writeCSR;
  wire                cpuClockingArea_rob_io_csrCtrl_ertn;
  wire                cpuClockingArea_rob_io_csrCtrl_normalException;
  wire                cpuClockingArea_rob_io_csrCtrl_tlbrException;
  wire       [31:0]   cpuClockingArea_rob_io_csrCtrl_epc;
  wire       [4:0]    cpuClockingArea_rob_io_csrCtrl_eROBIdx;
  wire       [5:0]    cpuClockingArea_rob_io_csrCtrl_eCode;
  wire       [0:0]    cpuClockingArea_rob_io_csrCtrl_eSubCode;
  wire                cpuClockingArea_rob_io_flush;
  wire       [31:0]   cpuClockingArea_rob_io_redirectPC;
  wire       [31:0]   cpuClockingArea_rob_io_commitROBEntries_0_pc;
  wire       [4:0]    cpuClockingArea_rob_io_commitROBEntries_0_ard;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_0_prd;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_0_pprd;
  wire       [3:0]    cpuClockingArea_rob_io_commitROBEntries_0_specialOp;
  wire                cpuClockingArea_rob_io_commitROBEntries_0_isComplete;
  wire       [31:0]   cpuClockingArea_rob_io_commitROBEntries_0_branchResult_targetPC;
  wire                cpuClockingArea_rob_io_commitROBEntries_0_branchResult_branchResult;
  wire                cpuClockingArea_rob_io_commitROBEntries_0_branchResult_predictFail;
  wire                cpuClockingArea_rob_io_commitROBEntries_0_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_0_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_rob_io_commitROBEntries_0_exceptionInfo_eSubCode;
  wire                cpuClockingArea_rob_io_commitROBEntries_0_valid;
  wire       [31:0]   cpuClockingArea_rob_io_commitROBEntries_1_pc;
  wire       [4:0]    cpuClockingArea_rob_io_commitROBEntries_1_ard;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_1_prd;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_1_pprd;
  wire       [3:0]    cpuClockingArea_rob_io_commitROBEntries_1_specialOp;
  wire                cpuClockingArea_rob_io_commitROBEntries_1_isComplete;
  wire       [31:0]   cpuClockingArea_rob_io_commitROBEntries_1_branchResult_targetPC;
  wire                cpuClockingArea_rob_io_commitROBEntries_1_branchResult_branchResult;
  wire                cpuClockingArea_rob_io_commitROBEntries_1_branchResult_predictFail;
  wire                cpuClockingArea_rob_io_commitROBEntries_1_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_1_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_rob_io_commitROBEntries_1_exceptionInfo_eSubCode;
  wire                cpuClockingArea_rob_io_commitROBEntries_1_valid;
  wire       [31:0]   cpuClockingArea_rob_io_commitROBEntries_2_pc;
  wire       [4:0]    cpuClockingArea_rob_io_commitROBEntries_2_ard;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_2_prd;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_2_pprd;
  wire       [3:0]    cpuClockingArea_rob_io_commitROBEntries_2_specialOp;
  wire                cpuClockingArea_rob_io_commitROBEntries_2_isComplete;
  wire       [31:0]   cpuClockingArea_rob_io_commitROBEntries_2_branchResult_targetPC;
  wire                cpuClockingArea_rob_io_commitROBEntries_2_branchResult_branchResult;
  wire                cpuClockingArea_rob_io_commitROBEntries_2_branchResult_predictFail;
  wire                cpuClockingArea_rob_io_commitROBEntries_2_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_2_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_rob_io_commitROBEntries_2_exceptionInfo_eSubCode;
  wire                cpuClockingArea_rob_io_commitROBEntries_2_valid;
  wire       [31:0]   cpuClockingArea_rob_io_commitROBEntries_3_pc;
  wire       [4:0]    cpuClockingArea_rob_io_commitROBEntries_3_ard;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_3_prd;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_3_pprd;
  wire       [3:0]    cpuClockingArea_rob_io_commitROBEntries_3_specialOp;
  wire                cpuClockingArea_rob_io_commitROBEntries_3_isComplete;
  wire       [31:0]   cpuClockingArea_rob_io_commitROBEntries_3_branchResult_targetPC;
  wire                cpuClockingArea_rob_io_commitROBEntries_3_branchResult_branchResult;
  wire                cpuClockingArea_rob_io_commitROBEntries_3_branchResult_predictFail;
  wire                cpuClockingArea_rob_io_commitROBEntries_3_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_3_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_rob_io_commitROBEntries_3_exceptionInfo_eSubCode;
  wire                cpuClockingArea_rob_io_commitROBEntries_3_valid;
  wire       [31:0]   cpuClockingArea_rob_io_commitROBEntries_4_pc;
  wire       [4:0]    cpuClockingArea_rob_io_commitROBEntries_4_ard;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_4_prd;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_4_pprd;
  wire       [3:0]    cpuClockingArea_rob_io_commitROBEntries_4_specialOp;
  wire                cpuClockingArea_rob_io_commitROBEntries_4_isComplete;
  wire       [31:0]   cpuClockingArea_rob_io_commitROBEntries_4_branchResult_targetPC;
  wire                cpuClockingArea_rob_io_commitROBEntries_4_branchResult_branchResult;
  wire                cpuClockingArea_rob_io_commitROBEntries_4_branchResult_predictFail;
  wire                cpuClockingArea_rob_io_commitROBEntries_4_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_rob_io_commitROBEntries_4_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_rob_io_commitROBEntries_4_exceptionInfo_eSubCode;
  wire                cpuClockingArea_rob_io_commitROBEntries_4_valid;
  wire                cpuClockingArea_csr_io_interrupt;
  wire       [1:0]    cpuClockingArea_csr__zz_when_Cache_l83;
  wire       [31:0]   cpuClockingArea_csr_io_counter_id;
  wire       [63:0]   cpuClockingArea_csr_io_counter_value;
  wire       [31:0]   cpuClockingArea_csr_io_swRead_value;
  wire       [31:0]   cpuClockingArea_csr_io_llBitComm_actualAddr;
  wire                cpuClockingArea_csr__zz_scMatchHit;
  wire       [9:0]    cpuClockingArea_csr_io_tlbCSRInfo_asid;
  wire       [1:0]    cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_plv;
  wire                cpuClockingArea_csr__zz_when_TLB_l177;
  wire                cpuClockingArea_csr__zz_when_TLB_l177_1;
  wire       [1:0]    cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_mat;
  wire       [1:0]    cpuClockingArea_csr__zz_io_dCacheReq_pageInfo_mat;
  wire                cpuClockingArea_csr__zz_when_TLB_l178;
  wire                cpuClockingArea_csr__zz_when_TLB_l178_1;
  wire       [1:0]    cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_mat_1;
  wire       [2:0]    cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_ppn;
  wire       [2:0]    cpuClockingArea_csr__zz_when_TLB_l178_2;
  wire                cpuClockingArea_csr__zz_when_TLB_l185;
  wire                cpuClockingArea_csr__zz_when_TLB_l185_1;
  wire       [1:0]    cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_mat_2;
  wire       [2:0]    cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_ppn_1;
  wire       [2:0]    cpuClockingArea_csr__zz_when_TLB_l185_2;
  wire       [5:0]    cpuClockingArea_csr__zz_entryToFill_e;
  wire       [1:0]    cpuClockingArea_csr__zz_io_csrWrite_asid;
  wire       [21:0]   cpuClockingArea_csr__zz_io_swRead_value;
  wire       [5:0]    cpuClockingArea_csr__zz_entryToFill_ps;
  wire                cpuClockingArea_csr__zz_io_swRead_value_1;
  wire                cpuClockingArea_csr__zz_entryToFill_e_1;
  wire       [18:0]   cpuClockingArea_csr__zz_entryToFill_vppn;
  wire                cpuClockingArea_csr__zz_entryToFill_pp0_v;
  wire                cpuClockingArea_csr__zz_entryToFill_pp0_d;
  wire       [1:0]    cpuClockingArea_csr__zz_entryToFill_pp0_plv;
  wire       [1:0]    cpuClockingArea_csr__zz_entryToFill_pp0_mat;
  wire                cpuClockingArea_csr__zz_entryToFill_g;
  wire       [19:0]   cpuClockingArea_csr__zz_entryToFill_pp0_ppn;
  wire                cpuClockingArea_csr__zz_entryToFill_pp1_v;
  wire                cpuClockingArea_csr__zz_entryToFill_pp1_d;
  wire       [1:0]    cpuClockingArea_csr__zz_entryToFill_pp1_plv;
  wire       [1:0]    cpuClockingArea_csr__zz_entryToFill_pp1_mat;
  wire                cpuClockingArea_csr__zz_entryToFill_g_1;
  wire       [19:0]   cpuClockingArea_csr__zz_entryToFill_pp1_ppn;
  wire       [31:0]   cpuClockingArea_csr_io_ctrl_era;
  wire       [31:0]   cpuClockingArea_csr_io_ctrl_eentry;
  wire       [31:0]   cpuClockingArea_csr_io_ctrl_tlbrentry;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_crmd;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_prmd;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_ecfg;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_estat;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_era;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_badv;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_eentry;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_tlbidx;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_tlbehi;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_tlbelo0;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_tlbelo1;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_asid;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_pgdl;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_pgdh;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_save0;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_save1;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_save2;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_save3;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_tid;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_tcfg;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_tval;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_ticlr;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_llbctl;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_tlbrentry;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_dmw0;
  wire       [31:0]   cpuClockingArea_csr_io_diffCSRBundle_dmw1;
  wire       [1:0]    cpuClockingArea_areaFlushReset_instQueue_io_in_allowMask;
  wire       [1:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_availMask;
  wire       [31:0]   cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_inst;
  wire       [31:0]   cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_branchInfo_predictPC;
  wire                cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_branchInfo_predictResult;
  wire                cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_pc;
  wire       [31:0]   cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_inst;
  wire       [31:0]   cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_branchInfo_predictPC;
  wire                cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_branchInfo_predictResult;
  wire                cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_pc;
  wire       [2:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_fuType;
  wire       [4:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_ard;
  wire       [4:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_asrc_0;
  wire       [4:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_asrc_1;
  wire       [2:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_fuType;
  wire       [4:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_ard;
  wire       [4:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_asrc_0;
  wire       [4:0]    cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_asrc_1;
  wire       [1:0]    cpuClockingArea_areaFlushReset_dispatcher_io_input_allowMask;
  wire       [1:0]    cpuClockingArea_areaFlushReset_dispatcher_io_rob_allowMask;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_rob_pc_0;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_rob_pc_1;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_rob_ard_0;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_rob_ard_1;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_rob_prd_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_rob_prd_1;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_rob_pprd_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_rob_pprd_1;
  wire       [3:0]    cpuClockingArea_areaFlushReset_dispatcher_io_rob_specialOp_0;
  wire       [3:0]    cpuClockingArea_areaFlushReset_dispatcher_io_rob_specialOp_1;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_0_prd;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_0_ard;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_0_wen;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_1_prd;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_1_ard;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_1_wen;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_0_0_ard;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_0_1_ard;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_1_0_ard;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_1_1_ard;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_sratReadPPRD_0_ard;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_sratReadPPRD_1_ard;
  wire       [1:0]    cpuClockingArea_areaFlushReset_dispatcher_io_freelist_disPatchNum;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_branchInfo_predictPC;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_branchInfo_predictResult;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_prd;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_psrc_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_psrc_1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_imm;
  wire       [3:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_uop_aluOp;
  wire       [1:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_uop_bruOp;
  wire       [1:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_uop_cruOp;
  wire       [2:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_roop_aluROOp;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_srcReady_0;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_srcReady_1;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_branchInfo_predictPC;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_branchInfo_predictResult;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_prd;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_psrc_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_psrc_1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_imm;
  wire       [3:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_uop_aluOp;
  wire       [1:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_uop_bruOp;
  wire       [2:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_roop_aluROOp;
  wire       [1:0]    cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_roop_cruROOp;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_srcReady_0;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_srcReady_1;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_prd;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_psrc_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_psrc_1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_imm;
  wire       [1:0]    cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_uop_muluOp;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_srcReady_0;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_srcReady_1;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_prd;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_psrc_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_psrc_1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_imm;
  wire       [1:0]    cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_uop_divuOp;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_srcReady_0;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_srcReady_1;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_prd;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_psrc_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_psrc_1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_imm;
  wire       [3:0]    cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_uop_lsuOp;
  wire       [4:0]    cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_uop_lsuCoOp;
  wire       [0:0]    cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_roop_lsuROOp;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_srcReady_0;
  wire                cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_srcReady_1;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU0_io_input_ready;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU0_io_csrInQueue;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_branchInfo_predictPC;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_branchInfo_predictResult;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_prd;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_psrc_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_psrc_1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_imm;
  wire       [3:0]    cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_uop_aluOp;
  wire       [1:0]    cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_uop_bruOp;
  wire       [1:0]    cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_uop_cruOp;
  wire       [2:0]    cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_roop_aluROOp;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU0_io_wakeOut_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueALU0_io_wakeOut_payload;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU1_io_input_ready;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU1_io_csrInQueue;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_branchInfo_predictPC;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_branchInfo_predictResult;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_prd;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_psrc_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_psrc_1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_imm;
  wire       [3:0]    cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_uop_aluOp;
  wire       [1:0]    cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_uop_bruOp;
  wire       [2:0]    cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_roop_aluROOp;
  wire       [1:0]    cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_roop_cruROOp;
  wire                cpuClockingArea_areaFlushReset_issueQueueALU1_io_wakeOut_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueALU1_io_wakeOut_payload;
  wire                cpuClockingArea_areaFlushReset_issueQueueMULU_io_input_ready;
  wire                cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_prd;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_psrc_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_psrc_1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_imm;
  wire       [1:0]    cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_uop_muluOp;
  wire                cpuClockingArea_areaFlushReset_issueQueueDIVU_io_input_ready;
  wire                cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_prd;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_psrc_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_psrc_1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_imm;
  wire       [1:0]    cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_uop_divuOp;
  wire                cpuClockingArea_areaFlushReset_issueQueueLSU_io_input_ready;
  wire                cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_prd;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_psrc_0;
  wire       [5:0]    cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_psrc_1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_imm;
  wire       [3:0]    cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_uop_lsuOp;
  wire       [4:0]    cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_uop_lsuCoOp;
  wire       [0:0]    cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_roop_lsuROOp;
  wire                cpuClockingArea_areaFlushReset_roALU0_io_cmd_ready;
  wire                cpuClockingArea_areaFlushReset_roALU0_io_toFU_valid;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src2;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src3;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src4;
  wire       [4:0]    cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_branchInfo_predictPC;
  wire                cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_branchInfo_predictResult;
  wire                cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_prd;
  wire       [3:0]    cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_uop_aluOp;
  wire       [1:0]    cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_uop_bruOp;
  wire       [1:0]    cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_uop_cruOp;
  wire                cpuClockingArea_areaFlushReset_roALU0_io_wakeOut_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roALU0_io_wakeOut_payload;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roALU0_io_prf_0_idx;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roALU0_io_prf_1_idx;
  wire       [13:0]   cpuClockingArea_areaFlushReset_roALU0_io_csr_address;
  wire                cpuClockingArea_areaFlushReset_roALU1_io_cmd_ready;
  wire                cpuClockingArea_areaFlushReset_roALU1_io_toFU_valid;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src2;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src3;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src4;
  wire       [4:0]    cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_branchInfo_predictPC;
  wire                cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_branchInfo_predictResult;
  wire                cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_prd;
  wire       [3:0]    cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_uop_aluOp;
  wire       [1:0]    cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_uop_bruOp;
  wire                cpuClockingArea_areaFlushReset_roALU1_io_wakeOut_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roALU1_io_wakeOut_payload;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roALU1_io_prf_0_idx;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roALU1_io_prf_1_idx;
  wire                cpuClockingArea_areaFlushReset_roMULU_io_cmd_ready;
  wire                cpuClockingArea_areaFlushReset_roMULU_io_toFU_valid;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_src1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_src2;
  wire       [4:0]    cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_prd;
  wire       [1:0]    cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_uop_muluOp;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roMULU_io_prf_0_idx;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roMULU_io_prf_1_idx;
  wire                cpuClockingArea_areaFlushReset_roDIVU_io_cmd_ready;
  wire                cpuClockingArea_areaFlushReset_roDIVU_io_toFU_valid;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_src1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_src2;
  wire       [4:0]    cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_prd;
  wire       [1:0]    cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_uop_divuOp;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roDIVU_io_prf_0_idx;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roDIVU_io_prf_1_idx;
  wire                cpuClockingArea_areaFlushReset_roLSU_io_cmd_ready;
  wire                cpuClockingArea_areaFlushReset_roLSU_io_toFU_valid;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_src1;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_src2;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_src3;
  wire       [4:0]    cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_exceptionInfo_eSubCode;
  wire       [31:0]   cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_pc;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_prd;
  wire       [3:0]    cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_uop_lsuOp;
  wire       [4:0]    cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_uop_lsuCoOp;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roLSU_io_prf_0_idx;
  wire       [5:0]    cpuClockingArea_areaFlushReset_roLSU_io_prf_1_idx;
  wire                cpuClockingArea_areaFlushReset_fuALU0_io_input_ready;
  wire                cpuClockingArea_areaFlushReset_fuALU0_io_output_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_data;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_prd;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_exceptionInfo_eSubCode;
  wire                cpuClockingArea_areaFlushReset_fuALU0_io_forward_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuALU0_io_forward_payload_idx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuALU0_io_forward_payload_payload;
  wire                cpuClockingArea_areaFlushReset_fuALU0_io_wakeOut_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuALU0_io_wakeOut_payload;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuALU0_io_csrWrite_value;
  wire       [13:0]   cpuClockingArea_areaFlushReset_fuALU0_io_csrWrite_address;
  wire                cpuClockingArea_areaFlushReset_fuALU0_io_csrWrite_wen;
  wire                cpuClockingArea_areaFlushReset_fuALU1_io_input_ready;
  wire                cpuClockingArea_areaFlushReset_fuALU1_io_output_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_data;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_prd;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_exceptionInfo_eSubCode;
  wire                cpuClockingArea_areaFlushReset_fuALU1_io_forward_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuALU1_io_forward_payload_idx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuALU1_io_forward_payload_payload;
  wire                cpuClockingArea_areaFlushReset_fuALU1_io_wakeOut_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuALU1_io_wakeOut_payload;
  wire                cpuClockingArea_areaFlushReset_fuMULU_io_input_ready;
  wire                cpuClockingArea_areaFlushReset_fuMULU_io_output_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_data;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_prd;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_exceptionInfo_eSubCode;
  wire                cpuClockingArea_areaFlushReset_fuMULU_io_forward_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuMULU_io_forward_payload_idx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuMULU_io_forward_payload_payload;
  wire                cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_0_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_0_payload;
  wire                cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_1_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_1_payload;
  wire                cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_2_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_2_payload;
  wire                cpuClockingArea_areaFlushReset_fuDIVU_io_input_ready;
  wire                cpuClockingArea_areaFlushReset_fuDIVU_io_output_valid;
  wire       [4:0]    cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_data;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_prd;
  wire       [31:0]   cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_exceptionInfo_eSubCode;
  wire                cpuClockingArea_areaFlushReset_commitALU0_io_input_ready;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitALU0_io_srat_prd;
  wire                cpuClockingArea_areaFlushReset_commitALU0_io_srat_wen;
  wire       [4:0]    cpuClockingArea_areaFlushReset_commitALU0_io_rob_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitALU0_io_rob_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_commitALU0_io_rob_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_commitALU0_io_rob_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_commitALU0_io_rob_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitALU0_io_rob_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_commitALU0_io_rob_exceptionInfo_eSubCode;
  wire                cpuClockingArea_areaFlushReset_commitALU0_io_rob_valid;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitALU0_io_prf_data;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitALU0_io_prf_idx;
  wire                cpuClockingArea_areaFlushReset_commitALU0_io_forward_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitALU0_io_forward_payload_idx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitALU0_io_forward_payload_payload;
  wire                cpuClockingArea_areaFlushReset_commitALU1_io_input_ready;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitALU1_io_srat_prd;
  wire                cpuClockingArea_areaFlushReset_commitALU1_io_srat_wen;
  wire       [4:0]    cpuClockingArea_areaFlushReset_commitALU1_io_rob_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitALU1_io_rob_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_commitALU1_io_rob_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_commitALU1_io_rob_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_commitALU1_io_rob_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitALU1_io_rob_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_commitALU1_io_rob_exceptionInfo_eSubCode;
  wire                cpuClockingArea_areaFlushReset_commitALU1_io_rob_valid;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitALU1_io_prf_data;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitALU1_io_prf_idx;
  wire                cpuClockingArea_areaFlushReset_commitALU1_io_forward_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitALU1_io_forward_payload_idx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitALU1_io_forward_payload_payload;
  wire                cpuClockingArea_areaFlushReset_commitMULU_io_input_ready;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitMULU_io_srat_prd;
  wire                cpuClockingArea_areaFlushReset_commitMULU_io_srat_wen;
  wire       [4:0]    cpuClockingArea_areaFlushReset_commitMULU_io_rob_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitMULU_io_rob_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_commitMULU_io_rob_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_commitMULU_io_rob_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_commitMULU_io_rob_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitMULU_io_rob_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_commitMULU_io_rob_exceptionInfo_eSubCode;
  wire                cpuClockingArea_areaFlushReset_commitMULU_io_rob_valid;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitMULU_io_prf_data;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitMULU_io_prf_idx;
  wire                cpuClockingArea_areaFlushReset_commitMULU_io_forward_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitMULU_io_forward_payload_idx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitMULU_io_forward_payload_payload;
  wire                cpuClockingArea_areaFlushReset_commitDIVU_io_input_ready;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitDIVU_io_srat_prd;
  wire                cpuClockingArea_areaFlushReset_commitDIVU_io_srat_wen;
  wire       [4:0]    cpuClockingArea_areaFlushReset_commitDIVU_io_rob_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitDIVU_io_rob_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_commitDIVU_io_rob_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_commitDIVU_io_rob_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_commitDIVU_io_rob_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitDIVU_io_rob_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_commitDIVU_io_rob_exceptionInfo_eSubCode;
  wire                cpuClockingArea_areaFlushReset_commitDIVU_io_rob_valid;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitDIVU_io_prf_data;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitDIVU_io_prf_idx;
  wire                cpuClockingArea_areaFlushReset_commitDIVU_io_forward_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitDIVU_io_forward_payload_idx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitDIVU_io_forward_payload_payload;
  wire                cpuClockingArea_areaFlushReset_commitLSU_io_input_ready;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitLSU_io_srat_prd;
  wire                cpuClockingArea_areaFlushReset_commitLSU_io_srat_wen;
  wire       [4:0]    cpuClockingArea_areaFlushReset_commitLSU_io_rob_robIdx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitLSU_io_rob_branchResult_targetPC;
  wire                cpuClockingArea_areaFlushReset_commitLSU_io_rob_branchResult_branchResult;
  wire                cpuClockingArea_areaFlushReset_commitLSU_io_rob_branchResult_predictFail;
  wire                cpuClockingArea_areaFlushReset_commitLSU_io_rob_exceptionInfo_exception;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitLSU_io_rob_exceptionInfo_eCode;
  wire       [0:0]    cpuClockingArea_areaFlushReset_commitLSU_io_rob_exceptionInfo_eSubCode;
  wire                cpuClockingArea_areaFlushReset_commitLSU_io_rob_valid;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitLSU_io_prf_data;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitLSU_io_prf_idx;
  wire                cpuClockingArea_areaFlushReset_commitLSU_io_forward_valid;
  wire       [5:0]    cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_idx;
  wire       [31:0]   cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_payload;
  reg        [31:0]   _zz_DaRAT_val_1;
  wire       [5:0]    _zz_DaRAT_val_1_1;
  reg        [31:0]   _zz_DaRAT_val_2;
  wire       [5:0]    _zz_DaRAT_val_2_1;
  reg        [31:0]   _zz_DaRAT_val_3;
  wire       [5:0]    _zz_DaRAT_val_3_1;
  reg        [31:0]   _zz_DaRAT_val_4;
  wire       [5:0]    _zz_DaRAT_val_4_1;
  reg        [31:0]   _zz_DaRAT_val_5;
  wire       [5:0]    _zz_DaRAT_val_5_1;
  reg        [31:0]   _zz_DaRAT_val_6;
  wire       [5:0]    _zz_DaRAT_val_6_1;
  reg        [31:0]   _zz_DaRAT_val_7;
  wire       [5:0]    _zz_DaRAT_val_7_1;
  reg        [31:0]   _zz_DaRAT_val_8;
  wire       [5:0]    _zz_DaRAT_val_8_1;
  reg        [31:0]   _zz_DaRAT_val_9;
  wire       [5:0]    _zz_DaRAT_val_9_1;
  reg        [31:0]   _zz_DaRAT_val_10;
  wire       [5:0]    _zz_DaRAT_val_10_1;
  reg        [31:0]   _zz_DaRAT_val_11;
  wire       [5:0]    _zz_DaRAT_val_11_1;
  reg        [31:0]   _zz_DaRAT_val_12;
  wire       [5:0]    _zz_DaRAT_val_12_1;
  reg        [31:0]   _zz_DaRAT_val_13;
  wire       [5:0]    _zz_DaRAT_val_13_1;
  reg        [31:0]   _zz_DaRAT_val_14;
  wire       [5:0]    _zz_DaRAT_val_14_1;
  reg        [31:0]   _zz_DaRAT_val_15;
  wire       [5:0]    _zz_DaRAT_val_15_1;
  reg        [31:0]   _zz_DaRAT_val_16;
  wire       [5:0]    _zz_DaRAT_val_16_1;
  reg        [31:0]   _zz_DaRAT_val_17;
  wire       [5:0]    _zz_DaRAT_val_17_1;
  reg        [31:0]   _zz_DaRAT_val_18;
  wire       [5:0]    _zz_DaRAT_val_18_1;
  reg        [31:0]   _zz_DaRAT_val_19;
  wire       [5:0]    _zz_DaRAT_val_19_1;
  reg        [31:0]   _zz_DaRAT_val_20;
  wire       [5:0]    _zz_DaRAT_val_20_1;
  reg        [31:0]   _zz_DaRAT_val_21;
  wire       [5:0]    _zz_DaRAT_val_21_1;
  reg        [31:0]   _zz_DaRAT_val_22;
  wire       [5:0]    _zz_DaRAT_val_22_1;
  reg        [31:0]   _zz_DaRAT_val_23;
  wire       [5:0]    _zz_DaRAT_val_23_1;
  reg        [31:0]   _zz_DaRAT_val_24;
  wire       [5:0]    _zz_DaRAT_val_24_1;
  reg        [31:0]   _zz_DaRAT_val_25;
  wire       [5:0]    _zz_DaRAT_val_25_1;
  reg        [31:0]   _zz_DaRAT_val_26;
  wire       [5:0]    _zz_DaRAT_val_26_1;
  reg        [31:0]   _zz_DaRAT_val_27;
  wire       [5:0]    _zz_DaRAT_val_27_1;
  reg        [31:0]   _zz_DaRAT_val_28;
  wire       [5:0]    _zz_DaRAT_val_28_1;
  reg        [31:0]   _zz_DaRAT_val_29;
  wire       [5:0]    _zz_DaRAT_val_29_1;
  reg        [31:0]   _zz_DaRAT_val_30;
  wire       [5:0]    _zz_DaRAT_val_30_1;
  reg        [31:0]   _zz_DaRAT_val_31;
  wire       [5:0]    _zz_DaRAT_val_31_1;
  wire       [31:0]   _zz_DifftestBundle_DifftestInstrCommitPC_0;
  wire       [31:0]   _zz_DifftestBundle_DifftestInstrCommitPC_1;
  wire       [31:0]   _zz_DifftestBundle_DifftestInstrCommitPC_2;
  wire       [31:0]   _zz_DifftestBundle_DifftestInstrCommitPC_3;
  wire       [31:0]   _zz_DifftestBundle_DifftestInstrCommitPC_4;
  wire       [1:0]    _zz_DifftestBundle_DifftestTlbFillIndex_4;
  wire       [31:0]   _zz_DifftestBundle_DifftestCount_1;
  wire       [31:0]   _zz_DifftestBundle_DifftestWdata_0;
  wire       [31:0]   _zz_DifftestBundle_DifftestWdata_1;
  wire       [31:0]   _zz_DifftestBundle_DifftestWdata_2;
  wire       [31:0]   _zz_DifftestBundle_DifftestWdata_3;
  wire       [31:0]   _zz_DifftestBundle_DifftestWdata_4;
  wire       [31:0]   _zz_DifftestBundle_DifftestExcpEventEPC;
  wire                cpuClockingArea_areaFlushReset_newReset;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_ready;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_branchInfo_predictPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_branchInfo_predictResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_pc;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_prd;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_psrc_0;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_psrc_1;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_imm;
  wire       [3:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp;
  wire       [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_bruOp;
  wire       [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_cruOp;
  wire       [2:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rValid;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_branchInfo_predictPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_branchInfo_predictResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_exceptionInfo_eSubCode;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_pc;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_prd;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_psrc_0;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_psrc_1;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_imm;
  reg        [3:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp;
  reg        [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_bruOp;
  reg        [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_cruOp;
  reg        [2:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp;
  wire                when_Stream_l369;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_ready;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_branchInfo_predictPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_branchInfo_predictResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_pc;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_prd;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_psrc_0;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_psrc_1;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_imm;
  wire       [3:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp;
  wire       [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_bruOp;
  wire       [2:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp;
  wire       [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_cruROOp;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rValid;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_branchInfo_predictPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_branchInfo_predictResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_exceptionInfo_eSubCode;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_pc;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_prd;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_psrc_0;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_psrc_1;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_imm;
  reg        [3:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp;
  reg        [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_bruOp;
  reg        [2:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp;
  reg        [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_cruROOp;
  wire                when_Stream_l369_1;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_ready;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_branchResult_targetPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_branchResult_branchResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_branchResult_predictFail;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_pc;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_prd;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_psrc_0;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_psrc_1;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_imm;
  wire       [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_uop_muluOp;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rValid;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_branchResult_targetPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_branchResult_branchResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_branchResult_predictFail;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_exceptionInfo_eSubCode;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_pc;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_prd;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_psrc_0;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_psrc_1;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_imm;
  reg        [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_uop_muluOp;
  wire                when_Stream_l369_2;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_ready;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_branchResult_targetPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_branchResult_branchResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_branchResult_predictFail;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_pc;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_prd;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_psrc_0;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_psrc_1;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_imm;
  wire       [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_uop_divuOp;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rValid;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_branchResult_targetPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_branchResult_branchResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_branchResult_predictFail;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_exceptionInfo_eSubCode;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_pc;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_prd;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_psrc_0;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_psrc_1;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_imm;
  reg        [1:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_uop_divuOp;
  wire                when_Stream_l369_3;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_ready;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_branchResult_targetPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_branchResult_branchResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_branchResult_predictFail;
  wire                toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_pc;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_prd;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_psrc_0;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_psrc_1;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_imm;
  wire       [3:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuCoOp;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_roop_lsuROOp;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rValid;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_branchResult_targetPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_branchResult_branchResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_branchResult_predictFail;
  reg                 toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_exceptionInfo_eSubCode;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_pc;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_prd;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_psrc_0;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_psrc_1;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_imm;
  reg        [3:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuCoOp;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_roop_lsuROOp;
  wire                when_Stream_l369_4;
  wire                toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_ready;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src1;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src2;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src3;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src4;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_branchInfo_predictPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_branchInfo_predictResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_pc;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_prd;
  wire       [3:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp;
  wire       [1:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_bruOp;
  wire       [1:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_cruOp;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rValid;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src1;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src2;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src3;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src4;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_branchInfo_predictPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_branchInfo_predictResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_exceptionInfo_eSubCode;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_pc;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_prd;
  reg        [3:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp;
  reg        [1:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_bruOp;
  reg        [1:0]    toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_cruOp;
  wire                when_Stream_l369_5;
  wire                toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_ready;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src1;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src2;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src3;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src4;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_branchInfo_predictPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_branchInfo_predictResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_pc;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_prd;
  wire       [3:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp;
  wire       [1:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_bruOp;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rValid;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src1;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src2;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src3;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src4;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_branchInfo_predictPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_branchInfo_predictResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_exceptionInfo_eSubCode;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_pc;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_prd;
  reg        [3:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp;
  reg        [1:0]    toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_bruOp;
  wire                when_Stream_l369_6;
  wire                toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_ready;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_src1;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_src2;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_branchResult_targetPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_branchResult_branchResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_branchResult_predictFail;
  wire                toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_pc;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_prd;
  wire       [1:0]    toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_uop_muluOp;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rValid;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_src1;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_src2;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_branchResult_targetPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_branchResult_branchResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_branchResult_predictFail;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_exceptionInfo_eSubCode;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_pc;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_prd;
  reg        [1:0]    toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_uop_muluOp;
  wire                when_Stream_l369_7;
  wire                toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_ready;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_src1;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_src2;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_branchResult_targetPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_branchResult_branchResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_branchResult_predictFail;
  wire                toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_pc;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_prd;
  wire       [1:0]    toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_uop_divuOp;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rValid;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_src1;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_src2;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_branchResult_targetPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_branchResult_branchResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_branchResult_predictFail;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_exceptionInfo_eSubCode;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_pc;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_prd;
  reg        [1:0]    toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_uop_divuOp;
  wire                when_Stream_l369_8;
  wire                toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_ready;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_src1;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_src2;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_src3;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_branchResult_targetPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_branchResult_branchResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_branchResult_predictFail;
  wire                toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_pc;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_prd;
  wire       [3:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuCoOp;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rValid;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_src1;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_src2;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_src3;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_branchResult_targetPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_branchResult_branchResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_branchResult_predictFail;
  reg                 toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_exceptionInfo_eSubCode;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_pc;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_prd;
  reg        [3:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuCoOp;
  wire                when_Stream_l369_9;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_ready;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_data;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_prd;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_branchResult_targetPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_branchResult_branchResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_branchResult_predictFail;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_exceptionInfo_eSubCode;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rValid;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_data;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_prd;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_branchResult_targetPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_branchResult_branchResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_branchResult_predictFail;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_exceptionInfo_eSubCode;
  wire                when_Stream_l369_10;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_ready;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_data;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_prd;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_branchResult_targetPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_branchResult_branchResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_branchResult_predictFail;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_exceptionInfo_eSubCode;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rValid;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_data;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_prd;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_branchResult_targetPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_branchResult_branchResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_branchResult_predictFail;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_exceptionInfo_eSubCode;
  wire                when_Stream_l369_11;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_ready;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_data;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_prd;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_branchResult_targetPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_branchResult_branchResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_branchResult_predictFail;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_exceptionInfo_eSubCode;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rValid;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_data;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_prd;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_branchResult_targetPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_branchResult_branchResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_branchResult_predictFail;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_exceptionInfo_eSubCode;
  wire                when_Stream_l369_12;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_ready;
  wire       [4:0]    toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_data;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_prd;
  wire       [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_branchResult_targetPC;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_branchResult_branchResult;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_branchResult_predictFail;
  wire                toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_exceptionInfo_eSubCode;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rValid;
  reg        [4:0]    toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_data;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_prd;
  reg        [31:0]   toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_branchResult_targetPC;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_branchResult_branchResult;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_branchResult_predictFail;
  reg                 toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_exceptionInfo_eSubCode;
  wire                when_Stream_l369_13;
  wire                toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_valid;
  wire                toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_ready;
  wire       [4:0]    toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_robIdx;
  wire       [31:0]   toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_data;
  wire       [5:0]    toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_prd;
  wire       [31:0]   toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_branchResult_targetPC;
  wire                toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_branchResult_branchResult;
  wire                toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_branchResult_predictFail;
  wire                toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_exceptionInfo_eSubCode;
  reg                 toplevel_cpuClockingArea_fuLSU_io_output_rValid;
  reg        [4:0]    toplevel_cpuClockingArea_fuLSU_io_output_rData_robIdx;
  reg        [31:0]   toplevel_cpuClockingArea_fuLSU_io_output_rData_data;
  reg        [5:0]    toplevel_cpuClockingArea_fuLSU_io_output_rData_prd;
  reg        [31:0]   toplevel_cpuClockingArea_fuLSU_io_output_rData_branchResult_targetPC;
  reg                 toplevel_cpuClockingArea_fuLSU_io_output_rData_branchResult_branchResult;
  reg                 toplevel_cpuClockingArea_fuLSU_io_output_rData_branchResult_predictFail;
  reg                 toplevel_cpuClockingArea_fuLSU_io_output_rData_exceptionInfo_exception;
  reg        [5:0]    toplevel_cpuClockingArea_fuLSU_io_output_rData_exceptionInfo_eCode;
  reg        [0:0]    toplevel_cpuClockingArea_fuLSU_io_output_rData_exceptionInfo_eSubCode;
  wire                when_Stream_l369_14;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_0_2;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_1_2;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_2_2;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_3_2;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_4_2;
  reg                 _zz_DifftestDelayBundle_DifftestInstrCommitValid_0_2;
  reg                 _zz_DifftestDelayBundle_DifftestInstrCommitValid_1_2;
  reg                 _zz_DifftestDelayBundle_DifftestInstrCommitValid_2_2;
  reg                 _zz_DifftestDelayBundle_DifftestInstrCommitValid_3_2;
  reg                 _zz_DifftestDelayBundle_DifftestInstrCommitValid_4_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_0_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_1_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_2_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_3_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestInstrCommitPC_4_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_0_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_1_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_2_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_3_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestInstrCommitInstr_4_2;
  reg                 _zz_DifftestDelayBundle_DifftestSkip_0_2;
  reg                 _zz_DifftestDelayBundle_DifftestSkip_1_2;
  reg                 _zz_DifftestDelayBundle_DifftestSkip_2_2;
  reg                 _zz_DifftestDelayBundle_DifftestSkip_3_2;
  reg                 _zz_DifftestDelayBundle_DifftestSkip_4_2;
  reg                 _zz_DifftestDelayBundle_DifftestIsTlbFill_0_2;
  reg                 _zz_DifftestDelayBundle_DifftestIsTlbFill_1_2;
  reg                 _zz_DifftestDelayBundle_DifftestIsTlbFill_2_2;
  reg                 _zz_DifftestDelayBundle_DifftestIsTlbFill_3_2;
  reg                 _zz_DifftestDelayBundle_DifftestIsTlbFill_4_2;
  reg        [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_0_2;
  reg        [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_1_2;
  reg        [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_2_2;
  reg        [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_3_2;
  reg        [4:0]    _zz_DifftestDelayBundle_DifftestTlbFillIndex_4_2;
  reg                 _zz_DifftestDelayBundle_DifftestIsCount_0_2;
  reg                 _zz_DifftestDelayBundle_DifftestIsCount_1_2;
  reg                 _zz_DifftestDelayBundle_DifftestIsCount_2_2;
  reg                 _zz_DifftestDelayBundle_DifftestIsCount_3_2;
  reg                 _zz_DifftestDelayBundle_DifftestIsCount_4_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestCount_0_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestCount_1_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestCount_2_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestCount_3_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestCount_4_2;
  reg                 _zz_DifftestDelayBundle_DifftestWen_0_2;
  reg                 _zz_DifftestDelayBundle_DifftestWen_1_2;
  reg                 _zz_DifftestDelayBundle_DifftestWen_2_2;
  reg                 _zz_DifftestDelayBundle_DifftestWen_3_2;
  reg                 _zz_DifftestDelayBundle_DifftestWen_4_2;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestWdest_0_2;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestWdest_1_2;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestWdest_2_2;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestWdest_3_2;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestWdest_4_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestWdata_0_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestWdata_1_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestWdata_2_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestWdata_3_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestWdata_4_2;
  reg                 _zz_DifftestDelayBundle_DifftestCsrRstat_0_2;
  reg                 _zz_DifftestDelayBundle_DifftestCsrRstat_1_2;
  reg                 _zz_DifftestDelayBundle_DifftestCsrRstat_2_2;
  reg                 _zz_DifftestDelayBundle_DifftestCsrRstat_3_2;
  reg                 _zz_DifftestDelayBundle_DifftestCsrRstat_4_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_0_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_1_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_2_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_3_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestCsrData_4_2;
  reg                 _zz_DifftestDelayBundle_DifftestExcpEventExcpValid_2;
  reg                 _zz_DifftestDelayBundle_DifftestExcpEventEret_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestExcpEventIntrNO_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestExcpEventCause_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestExcpEventEPC_2;
  reg        [31:0]   _zz_DifftestDelayBundle_DifftestExcpEventInst_2;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestStoreEventValid_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestStoreEventPAddr_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestStoreEventVAddr_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestStoreEventData_2;
  reg        [7:0]    _zz_DifftestDelayBundle_DifftestLoadEventValid_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestLoadEventPAddr_2;
  reg        [63:0]   _zz_DifftestDelayBundle_DifftestLoadEventVAddr_2;
  `ifndef SYNTHESIS
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_bruOp_string;
  reg [31:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_cruOp_string;
  reg [55:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_bruOp_string;
  reg [31:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_cruOp_string;
  reg [55:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_bruOp_string;
  reg [55:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp_string;
  reg [15:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_cruROOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_bruOp_string;
  reg [55:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp_string;
  reg [15:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_cruROOp_string;
  reg [47:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_uop_muluOp_string;
  reg [47:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_uop_muluOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_uop_divuOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_uop_divuOp_string;
  reg [55:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string;
  reg [47:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_roop_lsuROOp_string;
  reg [55:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string;
  reg [47:0] toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_roop_lsuROOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_bruOp_string;
  reg [31:0] toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_cruOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_bruOp_string;
  reg [31:0] toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_cruOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_bruOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_bruOp_string;
  reg [47:0] toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_uop_muluOp_string;
  reg [47:0] toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_uop_muluOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_uop_divuOp_string;
  reg [39:0] toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_uop_divuOp_string;
  reg [55:0] toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string;
  reg [55:0] toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string;
  `endif


  assign _zz_DifftestBundle_DifftestInstrCommitPC_0 = cpuClockingArea_rob_io_commitROBEntries_0_pc;
  assign _zz_DifftestBundle_DifftestInstrCommitPC_1 = cpuClockingArea_rob_io_commitROBEntries_1_pc;
  assign _zz_DifftestBundle_DifftestInstrCommitPC_2 = cpuClockingArea_rob_io_commitROBEntries_2_pc;
  assign _zz_DifftestBundle_DifftestInstrCommitPC_3 = cpuClockingArea_rob_io_commitROBEntries_3_pc;
  assign _zz_DifftestBundle_DifftestInstrCommitPC_4 = cpuClockingArea_rob_io_commitROBEntries_4_pc;
  assign _zz_DifftestBundle_DifftestTlbFillIndex_4 = cpuClockingArea_memService_io_TLBCtrl_index;
  assign _zz_DifftestBundle_DifftestCount_1 = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_data;
  assign _zz_DifftestBundle_DifftestWdata_0 = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_data;
  assign _zz_DifftestBundle_DifftestWdata_1 = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_data;
  assign _zz_DifftestBundle_DifftestWdata_2 = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_data;
  assign _zz_DifftestBundle_DifftestWdata_3 = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_data;
  assign _zz_DifftestBundle_DifftestWdata_4 = toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_data;
  assign _zz_DifftestBundle_DifftestExcpEventEPC = cpuClockingArea_rob_io_csrCtrl_epc;
  assign _zz_DaRAT_val_1_1 = cpuClockingArea_aRAT_io_recoveryPort_1;
  assign _zz_DaRAT_val_2_1 = cpuClockingArea_aRAT_io_recoveryPort_2;
  assign _zz_DaRAT_val_3_1 = cpuClockingArea_aRAT_io_recoveryPort_3;
  assign _zz_DaRAT_val_4_1 = cpuClockingArea_aRAT_io_recoveryPort_4;
  assign _zz_DaRAT_val_5_1 = cpuClockingArea_aRAT_io_recoveryPort_5;
  assign _zz_DaRAT_val_6_1 = cpuClockingArea_aRAT_io_recoveryPort_6;
  assign _zz_DaRAT_val_7_1 = cpuClockingArea_aRAT_io_recoveryPort_7;
  assign _zz_DaRAT_val_8_1 = cpuClockingArea_aRAT_io_recoveryPort_8;
  assign _zz_DaRAT_val_9_1 = cpuClockingArea_aRAT_io_recoveryPort_9;
  assign _zz_DaRAT_val_10_1 = cpuClockingArea_aRAT_io_recoveryPort_10;
  assign _zz_DaRAT_val_11_1 = cpuClockingArea_aRAT_io_recoveryPort_11;
  assign _zz_DaRAT_val_12_1 = cpuClockingArea_aRAT_io_recoveryPort_12;
  assign _zz_DaRAT_val_13_1 = cpuClockingArea_aRAT_io_recoveryPort_13;
  assign _zz_DaRAT_val_14_1 = cpuClockingArea_aRAT_io_recoveryPort_14;
  assign _zz_DaRAT_val_15_1 = cpuClockingArea_aRAT_io_recoveryPort_15;
  assign _zz_DaRAT_val_16_1 = cpuClockingArea_aRAT_io_recoveryPort_16;
  assign _zz_DaRAT_val_17_1 = cpuClockingArea_aRAT_io_recoveryPort_17;
  assign _zz_DaRAT_val_18_1 = cpuClockingArea_aRAT_io_recoveryPort_18;
  assign _zz_DaRAT_val_19_1 = cpuClockingArea_aRAT_io_recoveryPort_19;
  assign _zz_DaRAT_val_20_1 = cpuClockingArea_aRAT_io_recoveryPort_20;
  assign _zz_DaRAT_val_21_1 = cpuClockingArea_aRAT_io_recoveryPort_21;
  assign _zz_DaRAT_val_22_1 = cpuClockingArea_aRAT_io_recoveryPort_22;
  assign _zz_DaRAT_val_23_1 = cpuClockingArea_aRAT_io_recoveryPort_23;
  assign _zz_DaRAT_val_24_1 = cpuClockingArea_aRAT_io_recoveryPort_24;
  assign _zz_DaRAT_val_25_1 = cpuClockingArea_aRAT_io_recoveryPort_25;
  assign _zz_DaRAT_val_26_1 = cpuClockingArea_aRAT_io_recoveryPort_26;
  assign _zz_DaRAT_val_27_1 = cpuClockingArea_aRAT_io_recoveryPort_27;
  assign _zz_DaRAT_val_28_1 = cpuClockingArea_aRAT_io_recoveryPort_28;
  assign _zz_DaRAT_val_29_1 = cpuClockingArea_aRAT_io_recoveryPort_29;
  assign _zz_DaRAT_val_30_1 = cpuClockingArea_aRAT_io_recoveryPort_30;
  assign _zz_DaRAT_val_31_1 = cpuClockingArea_aRAT_io_recoveryPort_31;
  AXIArbiter cpuClockingArea_arbiter (
    .io_out_arid       (cpuClockingArea_arbiter_io_out_arid[3:0]     ), //o
    .io_out_araddr     (cpuClockingArea_arbiter_io_out_araddr[31:0]  ), //o
    .io_out_arlen      (cpuClockingArea_arbiter_io_out_arlen[7:0]    ), //o
    .io_out_arsize     (cpuClockingArea_arbiter_io_out_arsize[2:0]   ), //o
    .io_out_arburst    (cpuClockingArea_arbiter_io_out_arburst[1:0]  ), //o
    .io_out_arlock     (cpuClockingArea_arbiter_io_out_arlock[1:0]   ), //o
    .io_out_arcache    (cpuClockingArea_arbiter_io_out_arcache[3:0]  ), //o
    .io_out_arprot     (cpuClockingArea_arbiter_io_out_arprot[2:0]   ), //o
    .io_out_arvalid    (cpuClockingArea_arbiter_io_out_arvalid       ), //o
    .io_out_arready    (arready                                      ), //i
    .io_out_rid        (rid[3:0]                                     ), //i
    .io_out_rdata      (rdata[31:0]                                  ), //i
    .io_out_rresp      (rresp[1:0]                                   ), //i
    .io_out_rlast      (rlast                                        ), //i
    .io_out_rvalid     (rvalid                                       ), //i
    .io_out_rready     (cpuClockingArea_arbiter_io_out_rready        ), //o
    .io_out_awid       (cpuClockingArea_arbiter_io_out_awid[3:0]     ), //o
    .io_out_awaddr     (cpuClockingArea_arbiter_io_out_awaddr[31:0]  ), //o
    .io_out_awlen      (cpuClockingArea_arbiter_io_out_awlen[7:0]    ), //o
    .io_out_awsize     (cpuClockingArea_arbiter_io_out_awsize[2:0]   ), //o
    .io_out_awburst    (cpuClockingArea_arbiter_io_out_awburst[1:0]  ), //o
    .io_out_awlock     (cpuClockingArea_arbiter_io_out_awlock[1:0]   ), //o
    .io_out_awcache    (cpuClockingArea_arbiter_io_out_awcache[3:0]  ), //o
    .io_out_awprot     (cpuClockingArea_arbiter_io_out_awprot[2:0]   ), //o
    .io_out_awvalid    (cpuClockingArea_arbiter_io_out_awvalid       ), //o
    .io_out_awready    (awready                                      ), //i
    .io_out_wid        (cpuClockingArea_arbiter_io_out_wid[3:0]      ), //o
    .io_out_wdata      (cpuClockingArea_arbiter_io_out_wdata[31:0]   ), //o
    .io_out_wstrb      (cpuClockingArea_arbiter_io_out_wstrb[3:0]    ), //o
    .io_out_wlast      (cpuClockingArea_arbiter_io_out_wlast         ), //o
    .io_out_wvalid     (cpuClockingArea_arbiter_io_out_wvalid        ), //o
    .io_out_wready     (wready                                       ), //i
    .io_out_bid        (bid[3:0]                                     ), //i
    .io_out_bresp      (bresp[1:0]                                   ), //i
    .io_out_bvalid     (bvalid                                       ), //i
    .io_out_bready     (cpuClockingArea_arbiter_io_out_bready        ), //o
    .io_iCache_arid    (cpuClockingArea_iCache_io_axi_arid[3:0]      ), //i
    .io_iCache_araddr  (cpuClockingArea_iCache_io_axi_araddr[31:0]   ), //i
    .io_iCache_arlen   (cpuClockingArea_iCache_io_axi_arlen[7:0]     ), //i
    .io_iCache_arsize  (cpuClockingArea_iCache_io_axi_arsize[2:0]    ), //i
    .io_iCache_arburst (cpuClockingArea_iCache_io_axi_arburst[1:0]   ), //i
    .io_iCache_arlock  (cpuClockingArea_iCache_io_axi_arlock[1:0]    ), //i
    .io_iCache_arcache (cpuClockingArea_iCache_io_axi_arcache[3:0]   ), //i
    .io_iCache_arprot  (cpuClockingArea_iCache_io_axi_arprot[2:0]    ), //i
    .io_iCache_arvalid (cpuClockingArea_iCache_io_axi_arvalid        ), //i
    .io_iCache_arready (cpuClockingArea_arbiter_io_iCache_arready    ), //o
    .io_iCache_rid     (cpuClockingArea_arbiter_io_iCache_rid[3:0]   ), //o
    .io_iCache_rdata   (cpuClockingArea_arbiter_io_iCache_rdata[31:0]), //o
    .io_iCache_rresp   (cpuClockingArea_arbiter_io_iCache_rresp[1:0] ), //o
    .io_iCache_rlast   (cpuClockingArea_arbiter_io_iCache_rlast      ), //o
    .io_iCache_rvalid  (cpuClockingArea_arbiter_io_iCache_rvalid     ), //o
    .io_iCache_rready  (cpuClockingArea_iCache_io_axi_rready         ), //i
    .io_dCache_arid    (cpuClockingArea_fuLSU_io_axi_arid[3:0]       ), //i
    .io_dCache_araddr  (cpuClockingArea_fuLSU_io_axi_araddr[31:0]    ), //i
    .io_dCache_arlen   (cpuClockingArea_fuLSU_io_axi_arlen[7:0]      ), //i
    .io_dCache_arsize  (cpuClockingArea_fuLSU_io_axi_arsize[2:0]     ), //i
    .io_dCache_arburst (cpuClockingArea_fuLSU_io_axi_arburst[1:0]    ), //i
    .io_dCache_arlock  (cpuClockingArea_fuLSU_io_axi_arlock[1:0]     ), //i
    .io_dCache_arcache (cpuClockingArea_fuLSU_io_axi_arcache[3:0]    ), //i
    .io_dCache_arprot  (cpuClockingArea_fuLSU_io_axi_arprot[2:0]     ), //i
    .io_dCache_arvalid (cpuClockingArea_fuLSU_io_axi_arvalid         ), //i
    .io_dCache_arready (cpuClockingArea_arbiter_io_dCache_arready    ), //o
    .io_dCache_rid     (cpuClockingArea_arbiter_io_dCache_rid[3:0]   ), //o
    .io_dCache_rdata   (cpuClockingArea_arbiter_io_dCache_rdata[31:0]), //o
    .io_dCache_rresp   (cpuClockingArea_arbiter_io_dCache_rresp[1:0] ), //o
    .io_dCache_rlast   (cpuClockingArea_arbiter_io_dCache_rlast      ), //o
    .io_dCache_rvalid  (cpuClockingArea_arbiter_io_dCache_rvalid     ), //o
    .io_dCache_rready  (cpuClockingArea_fuLSU_io_axi_rready          ), //i
    .io_dCache_awid    (cpuClockingArea_fuLSU_io_axi_awid[3:0]       ), //i
    .io_dCache_awaddr  (cpuClockingArea_fuLSU_io_axi_awaddr[31:0]    ), //i
    .io_dCache_awlen   (cpuClockingArea_fuLSU_io_axi_awlen[7:0]      ), //i
    .io_dCache_awsize  (cpuClockingArea_fuLSU_io_axi_awsize[2:0]     ), //i
    .io_dCache_awburst (cpuClockingArea_fuLSU_io_axi_awburst[1:0]    ), //i
    .io_dCache_awlock  (cpuClockingArea_fuLSU_io_axi_awlock[1:0]     ), //i
    .io_dCache_awcache (cpuClockingArea_fuLSU_io_axi_awcache[3:0]    ), //i
    .io_dCache_awprot  (cpuClockingArea_fuLSU_io_axi_awprot[2:0]     ), //i
    .io_dCache_awvalid (cpuClockingArea_fuLSU_io_axi_awvalid         ), //i
    .io_dCache_awready (cpuClockingArea_arbiter_io_dCache_awready    ), //o
    .io_dCache_wid     (cpuClockingArea_fuLSU_io_axi_wid[3:0]        ), //i
    .io_dCache_wdata   (cpuClockingArea_fuLSU_io_axi_wdata[31:0]     ), //i
    .io_dCache_wstrb   (cpuClockingArea_fuLSU_io_axi_wstrb[3:0]      ), //i
    .io_dCache_wlast   (cpuClockingArea_fuLSU_io_axi_wlast           ), //i
    .io_dCache_wvalid  (cpuClockingArea_fuLSU_io_axi_wvalid          ), //i
    .io_dCache_wready  (cpuClockingArea_arbiter_io_dCache_wready     ), //o
    .io_dCache_bid     (cpuClockingArea_arbiter_io_dCache_bid[3:0]   ), //o
    .io_dCache_bresp   (cpuClockingArea_arbiter_io_dCache_bresp[1:0] ), //o
    .io_dCache_bvalid  (cpuClockingArea_arbiter_io_dCache_bvalid     ), //o
    .io_dCache_bready  (cpuClockingArea_fuLSU_io_axi_bready          )  //i
  );
  TLB cpuClockingArea_tlb (
    .io_iCacheReq_hit                (cpuClockingArea_tlb_io_iCacheReq_hit                    ), //o
    .io_iCacheReq_pageInfo_ppn       (cpuClockingArea_tlb_io_iCacheReq_pageInfo_ppn[19:0]     ), //o
    .io_iCacheReq_pageInfo_plv       (cpuClockingArea_tlb_io_iCacheReq_pageInfo_plv[1:0]      ), //o
    .io_iCacheReq_pageInfo_mat       (cpuClockingArea_tlb_io_iCacheReq_pageInfo_mat[1:0]      ), //o
    .io_iCacheReq_pageInfo_d         (cpuClockingArea_tlb_io_iCacheReq_pageInfo_d             ), //o
    .io_iCacheReq_pageInfo_v         (cpuClockingArea_tlb_io_iCacheReq_pageInfo_v             ), //o
    .io_iCacheReq_virtPageNumber     (cpuClockingArea_iCache_io_tlb_virtPageNumber[19:0]      ), //i
    .io_dCacheReq_hit                (cpuClockingArea_tlb_io_dCacheReq_hit                    ), //o
    .io_dCacheReq_pageInfo_ppn       (cpuClockingArea_tlb_io_dCacheReq_pageInfo_ppn[19:0]     ), //o
    .io_dCacheReq_pageInfo_plv       (cpuClockingArea_tlb_io_dCacheReq_pageInfo_plv[1:0]      ), //o
    .io_dCacheReq_pageInfo_mat       (cpuClockingArea_tlb_io_dCacheReq_pageInfo_mat[1:0]      ), //o
    .io_dCacheReq_pageInfo_d         (cpuClockingArea_tlb_io_dCacheReq_pageInfo_d             ), //o
    .io_dCacheReq_pageInfo_v         (cpuClockingArea_tlb_io_dCacheReq_pageInfo_v             ), //o
    .io_dCacheReq_virtPageNumber     (cpuClockingArea_fuLSU_io_tlb_virtPageNumber[19:0]       ), //i
    .io_csrInfo_asid                 (cpuClockingArea_csr_io_tlbCSRInfo_asid[9:0]             ), //i
    ._zz_io_iCacheReq_pageInfo_plv   (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_plv[1:0]  ), //i
    ._zz_when_TLB_l177               (cpuClockingArea_csr__zz_when_TLB_l177                   ), //i
    ._zz_when_TLB_l177_1             (cpuClockingArea_csr__zz_when_TLB_l177_1                 ), //i
    ._zz_io_iCacheReq_pageInfo_mat   (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_mat[1:0]  ), //i
    ._zz_io_dCacheReq_pageInfo_mat   (cpuClockingArea_csr__zz_io_dCacheReq_pageInfo_mat[1:0]  ), //i
    ._zz_when_TLB_l178               (cpuClockingArea_csr__zz_when_TLB_l178                   ), //i
    ._zz_when_TLB_l178_1             (cpuClockingArea_csr__zz_when_TLB_l178_1                 ), //i
    ._zz_io_iCacheReq_pageInfo_mat_1 (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_mat_1[1:0]), //i
    ._zz_io_iCacheReq_pageInfo_ppn   (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_ppn[2:0]  ), //i
    ._zz_when_TLB_l178_2             (cpuClockingArea_csr__zz_when_TLB_l178_2[2:0]            ), //i
    ._zz_when_TLB_l185               (cpuClockingArea_csr__zz_when_TLB_l185                   ), //i
    ._zz_when_TLB_l185_1             (cpuClockingArea_csr__zz_when_TLB_l185_1                 ), //i
    ._zz_io_iCacheReq_pageInfo_mat_2 (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_mat_2[1:0]), //i
    ._zz_io_iCacheReq_pageInfo_ppn_1 (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_ppn_1[2:0]), //i
    ._zz_when_TLB_l185_2             (cpuClockingArea_csr__zz_when_TLB_l185_2[2:0]            ), //i
    ._zz_entryToFill_e               (cpuClockingArea_csr__zz_entryToFill_e[5:0]              ), //i
    ._zz_io_csrWrite_asid            (cpuClockingArea_csr__zz_io_csrWrite_asid[1:0]           ), //i
    ._zz_io_swRead_value             (cpuClockingArea_csr__zz_io_swRead_value[21:0]           ), //i
    ._zz_entryToFill_ps              (cpuClockingArea_csr__zz_entryToFill_ps[5:0]             ), //i
    ._zz_io_swRead_value_1           (cpuClockingArea_csr__zz_io_swRead_value_1               ), //i
    ._zz_entryToFill_e_1             (cpuClockingArea_csr__zz_entryToFill_e_1                 ), //i
    ._zz_entryToFill_vppn            (cpuClockingArea_csr__zz_entryToFill_vppn[18:0]          ), //i
    ._zz_entryToFill_pp0_v           (cpuClockingArea_csr__zz_entryToFill_pp0_v               ), //i
    ._zz_entryToFill_pp0_d           (cpuClockingArea_csr__zz_entryToFill_pp0_d               ), //i
    ._zz_entryToFill_pp0_plv         (cpuClockingArea_csr__zz_entryToFill_pp0_plv[1:0]        ), //i
    ._zz_entryToFill_pp0_mat         (cpuClockingArea_csr__zz_entryToFill_pp0_mat[1:0]        ), //i
    ._zz_entryToFill_g               (cpuClockingArea_csr__zz_entryToFill_g                   ), //i
    ._zz_entryToFill_pp0_ppn         (cpuClockingArea_csr__zz_entryToFill_pp0_ppn[19:0]       ), //i
    ._zz_entryToFill_pp1_v           (cpuClockingArea_csr__zz_entryToFill_pp1_v               ), //i
    ._zz_entryToFill_pp1_d           (cpuClockingArea_csr__zz_entryToFill_pp1_d               ), //i
    ._zz_entryToFill_pp1_plv         (cpuClockingArea_csr__zz_entryToFill_pp1_plv[1:0]        ), //i
    ._zz_entryToFill_pp1_mat         (cpuClockingArea_csr__zz_entryToFill_pp1_mat[1:0]        ), //i
    ._zz_entryToFill_g_1             (cpuClockingArea_csr__zz_entryToFill_g_1                 ), //i
    ._zz_entryToFill_pp1_ppn         (cpuClockingArea_csr__zz_entryToFill_pp1_ppn[19:0]       ), //i
    ._zz_io_swRead_value_2           (cpuClockingArea_tlb__zz_io_swRead_value_2[1:0]          ), //o
    ._zz_io_swRead_value_3           (cpuClockingArea_tlb__zz_io_swRead_value_3[21:0]         ), //o
    ._zz_io_swRead_value_4           (cpuClockingArea_tlb__zz_io_swRead_value_4[5:0]          ), //o
    ._zz_io_swRead_value_5           (cpuClockingArea_tlb__zz_io_swRead_value_5               ), //o
    ._zz_io_swRead_value_6           (cpuClockingArea_tlb__zz_io_swRead_value_6               ), //o
    ._zz_io_swRead_value_7           (cpuClockingArea_tlb__zz_io_swRead_value_7[12:0]         ), //o
    ._zz_io_swRead_value_8           (cpuClockingArea_tlb__zz_io_swRead_value_8[18:0]         ), //o
    ._zz_io_swRead_value_9           (cpuClockingArea_tlb__zz_io_swRead_value_9               ), //o
    ._zz_io_swRead_value_10          (cpuClockingArea_tlb__zz_io_swRead_value_10              ), //o
    ._zz_io_swRead_value_11          (cpuClockingArea_tlb__zz_io_swRead_value_11[1:0]         ), //o
    ._zz_io_swRead_value_12          (cpuClockingArea_tlb__zz_io_swRead_value_12[1:0]         ), //o
    ._zz_io_swRead_value_13          (cpuClockingArea_tlb__zz_io_swRead_value_13              ), //o
    ._zz_io_swRead_value_14          (cpuClockingArea_tlb__zz_io_swRead_value_14              ), //o
    ._zz_io_swRead_value_15          (cpuClockingArea_tlb__zz_io_swRead_value_15[19:0]        ), //o
    ._zz_io_swRead_value_16          (cpuClockingArea_tlb__zz_io_swRead_value_16[3:0]         ), //o
    ._zz_io_swRead_value_17          (cpuClockingArea_tlb__zz_io_swRead_value_17              ), //o
    ._zz_io_swRead_value_18          (cpuClockingArea_tlb__zz_io_swRead_value_18              ), //o
    ._zz_io_swRead_value_19          (cpuClockingArea_tlb__zz_io_swRead_value_19[1:0]         ), //o
    ._zz_io_swRead_value_20          (cpuClockingArea_tlb__zz_io_swRead_value_20[1:0]         ), //o
    ._zz_io_swRead_value_21          (cpuClockingArea_tlb__zz_io_swRead_value_21              ), //o
    ._zz_io_swRead_value_22          (cpuClockingArea_tlb__zz_io_swRead_value_22              ), //o
    ._zz_io_swRead_value_23          (cpuClockingArea_tlb__zz_io_swRead_value_23[19:0]        ), //o
    ._zz_io_swRead_value_24          (cpuClockingArea_tlb__zz_io_swRead_value_24[3:0]         ), //o
    .io_csrWrite_asid                (cpuClockingArea_tlb_io_csrWrite_asid[9:0]               ), //o
    .io_csrWrite_idxWen              (cpuClockingArea_tlb_io_csrWrite_idxWen                  ), //o
    .io_csrWrite_entryWen            (cpuClockingArea_tlb_io_csrWrite_entryWen                ), //o
    .io_ctrl_op                      (cpuClockingArea_memService_io_TLBCtrl_op[2:0]           ), //i
    .io_ctrl_invGlobal               (cpuClockingArea_memService_io_TLBCtrl_invGlobal         ), //i
    .io_ctrl_invLocal                (cpuClockingArea_memService_io_TLBCtrl_invLocal          ), //i
    .io_ctrl_invLocalVAMatch         (cpuClockingArea_memService_io_TLBCtrl_invLocalVAMatch   ), //i
    .io_ctrl_invLocalVANotMatch      (cpuClockingArea_memService_io_TLBCtrl_invLocalVANotMatch), //i
    .io_ctrl_index                   (cpuClockingArea_memService_io_TLBCtrl_index[1:0]        ), //i
    .io_ctrl_invVA                   (cpuClockingArea_memService_io_TLBCtrl_invVA[18:0]       ), //i
    .io_ctrl_asid                    (cpuClockingArea_memService_io_TLBCtrl_asid[9:0]         ), //i
    .aclk                            (aclk                                                    ), //i
    .aresetn                         (aresetn                                                 )  //i
  );
  MemService cpuClockingArea_memService (
    .io_input_valid                     (cpuClockingArea_fuLSU_io_specialOpBufferUpdate_valid                   ), //i
    .io_input_payload_uop_lsuOp         (cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_uop_lsuOp[3:0]  ), //i
    .io_input_payload_uop_lsuCoOp       (cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_uop_lsuCoOp[4:0]), //i
    .io_input_payload_vaddr             (cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_vaddr[31:0]     ), //i
    .io_input_payload_asid              (cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_asid[9:0]       ), //i
    .io_iCacheCtrl_busy                 (cpuClockingArea_iCache_io_ctrl_busy                                    ), //i
    .io_iCacheCtrl_stall                (cpuClockingArea_memService_io_iCacheCtrl_stall                         ), //o
    .io_iCacheCtrl_cacopVA              (cpuClockingArea_memService_io_iCacheCtrl_cacopVA[31:0]                 ), //o
    .io_iCacheCtrl_cacopStoreTag        (cpuClockingArea_memService_io_iCacheCtrl_cacopStoreTag                 ), //o
    .io_iCacheCtrl_cacopIndexInvalidate (cpuClockingArea_memService_io_iCacheCtrl_cacopIndexInvalidate          ), //o
    .io_iCacheCtrl_cacopHitInvalidate   (cpuClockingArea_memService_io_iCacheCtrl_cacopHitInvalidate            ), //o
    .io_dCacheCtrl_busy                 (cpuClockingArea_fuLSU_io_ctrl_busy                                     ), //i
    .io_dCacheCtrl_stall                (cpuClockingArea_memService_io_dCacheCtrl_stall                         ), //o
    .io_dCacheCtrl_cacopVA              (cpuClockingArea_memService_io_dCacheCtrl_cacopVA[31:0]                 ), //o
    .io_dCacheCtrl_cacopStoreTag        (cpuClockingArea_memService_io_dCacheCtrl_cacopStoreTag                 ), //o
    .io_dCacheCtrl_cacopIndexInvalidate (cpuClockingArea_memService_io_dCacheCtrl_cacopIndexInvalidate          ), //o
    .io_dCacheCtrl_cacopHitInvalidate   (cpuClockingArea_memService_io_dCacheCtrl_cacopHitInvalidate            ), //o
    .io_TLBCtrl_op                      (cpuClockingArea_memService_io_TLBCtrl_op[2:0]                          ), //o
    .io_TLBCtrl_invGlobal               (cpuClockingArea_memService_io_TLBCtrl_invGlobal                        ), //o
    .io_TLBCtrl_invLocal                (cpuClockingArea_memService_io_TLBCtrl_invLocal                         ), //o
    .io_TLBCtrl_invLocalVAMatch         (cpuClockingArea_memService_io_TLBCtrl_invLocalVAMatch                  ), //o
    .io_TLBCtrl_invLocalVANotMatch      (cpuClockingArea_memService_io_TLBCtrl_invLocalVANotMatch               ), //o
    .io_TLBCtrl_index                   (cpuClockingArea_memService_io_TLBCtrl_index[1:0]                       ), //o
    .io_TLBCtrl_invVA                   (cpuClockingArea_memService_io_TLBCtrl_invVA[18:0]                      ), //o
    .io_TLBCtrl_asid                    (cpuClockingArea_memService_io_TLBCtrl_asid[9:0]                        ), //o
    .io_flush                           (cpuClockingArea_rob_io_flush                                           ), //i
    .io_wake                            (cpuClockingArea_rob_io_wakeupMem                                       ), //i
    .aclk                               (aclk                                                                   ), //i
    .aresetn                            (aresetn                                                                )  //i
  );
  SRAT cpuClockingArea_sRAT (
    .io_writePort_0_ard         (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_0_ard[4:0]    ), //i
    .io_writePort_0_prd         (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_0_prd[5:0]    ), //i
    .io_writePort_0_wen         (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_0_wen         ), //i
    .io_writePort_1_ard         (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_1_ard[4:0]    ), //i
    .io_writePort_1_prd         (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_1_prd[5:0]    ), //i
    .io_writePort_1_wen         (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_1_wen         ), //i
    .io_updatePort_0_prd        (cpuClockingArea_areaFlushReset_commitALU0_io_srat_prd[5:0]           ), //i
    .io_updatePort_0_wen        (cpuClockingArea_areaFlushReset_commitALU0_io_srat_wen                ), //i
    .io_updatePort_1_prd        (cpuClockingArea_areaFlushReset_commitALU1_io_srat_prd[5:0]           ), //i
    .io_updatePort_1_wen        (cpuClockingArea_areaFlushReset_commitALU1_io_srat_wen                ), //i
    .io_updatePort_2_prd        (cpuClockingArea_areaFlushReset_commitMULU_io_srat_prd[5:0]           ), //i
    .io_updatePort_2_wen        (cpuClockingArea_areaFlushReset_commitMULU_io_srat_wen                ), //i
    .io_updatePort_3_prd        (cpuClockingArea_areaFlushReset_commitDIVU_io_srat_prd[5:0]           ), //i
    .io_updatePort_3_wen        (cpuClockingArea_areaFlushReset_commitDIVU_io_srat_wen                ), //i
    .io_updatePort_4_prd        (cpuClockingArea_areaFlushReset_commitLSU_io_srat_prd[5:0]            ), //i
    .io_updatePort_4_wen        (cpuClockingArea_areaFlushReset_commitLSU_io_srat_wen                 ), //i
    .io_srcReadPort_0_0_ard     (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_0_0_ard[4:0]), //i
    .io_srcReadPort_0_0_prd     (cpuClockingArea_sRAT_io_srcReadPort_0_0_prd[5:0]                     ), //o
    .io_srcReadPort_0_0_valid   (cpuClockingArea_sRAT_io_srcReadPort_0_0_valid                        ), //o
    .io_srcReadPort_0_1_ard     (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_0_1_ard[4:0]), //i
    .io_srcReadPort_0_1_prd     (cpuClockingArea_sRAT_io_srcReadPort_0_1_prd[5:0]                     ), //o
    .io_srcReadPort_0_1_valid   (cpuClockingArea_sRAT_io_srcReadPort_0_1_valid                        ), //o
    .io_srcReadPort_1_0_ard     (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_1_0_ard[4:0]), //i
    .io_srcReadPort_1_0_prd     (cpuClockingArea_sRAT_io_srcReadPort_1_0_prd[5:0]                     ), //o
    .io_srcReadPort_1_0_valid   (cpuClockingArea_sRAT_io_srcReadPort_1_0_valid                        ), //o
    .io_srcReadPort_1_1_ard     (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_1_1_ard[4:0]), //i
    .io_srcReadPort_1_1_prd     (cpuClockingArea_sRAT_io_srcReadPort_1_1_prd[5:0]                     ), //o
    .io_srcReadPort_1_1_valid   (cpuClockingArea_sRAT_io_srcReadPort_1_1_valid                        ), //o
    .io_prevPRDReadPort_0_ard   (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadPPRD_0_ard[4:0] ), //i
    .io_prevPRDReadPort_0_prd   (cpuClockingArea_sRAT_io_prevPRDReadPort_0_prd[5:0]                   ), //o
    .io_prevPRDReadPort_0_valid (cpuClockingArea_sRAT_io_prevPRDReadPort_0_valid                      ), //o
    .io_prevPRDReadPort_1_ard   (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadPPRD_1_ard[4:0] ), //i
    .io_prevPRDReadPort_1_prd   (cpuClockingArea_sRAT_io_prevPRDReadPort_1_prd[5:0]                   ), //o
    .io_prevPRDReadPort_1_valid (cpuClockingArea_sRAT_io_prevPRDReadPort_1_valid                      ), //o
    .io_delayedRecovery         (cpuClockingArea_rob_io_retireFreeList_delayedFlush                   ), //i
    .io_recoveryPort_0          (cpuClockingArea_aRAT_io_recoveryPort_0[5:0]                          ), //i
    .io_recoveryPort_1          (cpuClockingArea_aRAT_io_recoveryPort_1[5:0]                          ), //i
    .io_recoveryPort_2          (cpuClockingArea_aRAT_io_recoveryPort_2[5:0]                          ), //i
    .io_recoveryPort_3          (cpuClockingArea_aRAT_io_recoveryPort_3[5:0]                          ), //i
    .io_recoveryPort_4          (cpuClockingArea_aRAT_io_recoveryPort_4[5:0]                          ), //i
    .io_recoveryPort_5          (cpuClockingArea_aRAT_io_recoveryPort_5[5:0]                          ), //i
    .io_recoveryPort_6          (cpuClockingArea_aRAT_io_recoveryPort_6[5:0]                          ), //i
    .io_recoveryPort_7          (cpuClockingArea_aRAT_io_recoveryPort_7[5:0]                          ), //i
    .io_recoveryPort_8          (cpuClockingArea_aRAT_io_recoveryPort_8[5:0]                          ), //i
    .io_recoveryPort_9          (cpuClockingArea_aRAT_io_recoveryPort_9[5:0]                          ), //i
    .io_recoveryPort_10         (cpuClockingArea_aRAT_io_recoveryPort_10[5:0]                         ), //i
    .io_recoveryPort_11         (cpuClockingArea_aRAT_io_recoveryPort_11[5:0]                         ), //i
    .io_recoveryPort_12         (cpuClockingArea_aRAT_io_recoveryPort_12[5:0]                         ), //i
    .io_recoveryPort_13         (cpuClockingArea_aRAT_io_recoveryPort_13[5:0]                         ), //i
    .io_recoveryPort_14         (cpuClockingArea_aRAT_io_recoveryPort_14[5:0]                         ), //i
    .io_recoveryPort_15         (cpuClockingArea_aRAT_io_recoveryPort_15[5:0]                         ), //i
    .io_recoveryPort_16         (cpuClockingArea_aRAT_io_recoveryPort_16[5:0]                         ), //i
    .io_recoveryPort_17         (cpuClockingArea_aRAT_io_recoveryPort_17[5:0]                         ), //i
    .io_recoveryPort_18         (cpuClockingArea_aRAT_io_recoveryPort_18[5:0]                         ), //i
    .io_recoveryPort_19         (cpuClockingArea_aRAT_io_recoveryPort_19[5:0]                         ), //i
    .io_recoveryPort_20         (cpuClockingArea_aRAT_io_recoveryPort_20[5:0]                         ), //i
    .io_recoveryPort_21         (cpuClockingArea_aRAT_io_recoveryPort_21[5:0]                         ), //i
    .io_recoveryPort_22         (cpuClockingArea_aRAT_io_recoveryPort_22[5:0]                         ), //i
    .io_recoveryPort_23         (cpuClockingArea_aRAT_io_recoveryPort_23[5:0]                         ), //i
    .io_recoveryPort_24         (cpuClockingArea_aRAT_io_recoveryPort_24[5:0]                         ), //i
    .io_recoveryPort_25         (cpuClockingArea_aRAT_io_recoveryPort_25[5:0]                         ), //i
    .io_recoveryPort_26         (cpuClockingArea_aRAT_io_recoveryPort_26[5:0]                         ), //i
    .io_recoveryPort_27         (cpuClockingArea_aRAT_io_recoveryPort_27[5:0]                         ), //i
    .io_recoveryPort_28         (cpuClockingArea_aRAT_io_recoveryPort_28[5:0]                         ), //i
    .io_recoveryPort_29         (cpuClockingArea_aRAT_io_recoveryPort_29[5:0]                         ), //i
    .io_recoveryPort_30         (cpuClockingArea_aRAT_io_recoveryPort_30[5:0]                         ), //i
    .io_recoveryPort_31         (cpuClockingArea_aRAT_io_recoveryPort_31[5:0]                         ), //i
    .aclk                       (aclk                                                                 ), //i
    .aresetn                    (aresetn                                                              )  //i
  );
  ARAT cpuClockingArea_aRAT (
    .io_retirePort_0_ard (cpuClockingArea_rob_io_retireARAT_0_ard[4:0]), //i
    .io_retirePort_0_prd (cpuClockingArea_rob_io_retireARAT_0_prd[5:0]), //i
    .io_retirePort_0_wen (cpuClockingArea_rob_io_retireARAT_0_wen     ), //i
    .io_retirePort_1_ard (cpuClockingArea_rob_io_retireARAT_1_ard[4:0]), //i
    .io_retirePort_1_prd (cpuClockingArea_rob_io_retireARAT_1_prd[5:0]), //i
    .io_retirePort_1_wen (cpuClockingArea_rob_io_retireARAT_1_wen     ), //i
    .io_recoveryPort_0   (cpuClockingArea_aRAT_io_recoveryPort_0[5:0] ), //o
    .io_recoveryPort_1   (cpuClockingArea_aRAT_io_recoveryPort_1[5:0] ), //o
    .io_recoveryPort_2   (cpuClockingArea_aRAT_io_recoveryPort_2[5:0] ), //o
    .io_recoveryPort_3   (cpuClockingArea_aRAT_io_recoveryPort_3[5:0] ), //o
    .io_recoveryPort_4   (cpuClockingArea_aRAT_io_recoveryPort_4[5:0] ), //o
    .io_recoveryPort_5   (cpuClockingArea_aRAT_io_recoveryPort_5[5:0] ), //o
    .io_recoveryPort_6   (cpuClockingArea_aRAT_io_recoveryPort_6[5:0] ), //o
    .io_recoveryPort_7   (cpuClockingArea_aRAT_io_recoveryPort_7[5:0] ), //o
    .io_recoveryPort_8   (cpuClockingArea_aRAT_io_recoveryPort_8[5:0] ), //o
    .io_recoveryPort_9   (cpuClockingArea_aRAT_io_recoveryPort_9[5:0] ), //o
    .io_recoveryPort_10  (cpuClockingArea_aRAT_io_recoveryPort_10[5:0]), //o
    .io_recoveryPort_11  (cpuClockingArea_aRAT_io_recoveryPort_11[5:0]), //o
    .io_recoveryPort_12  (cpuClockingArea_aRAT_io_recoveryPort_12[5:0]), //o
    .io_recoveryPort_13  (cpuClockingArea_aRAT_io_recoveryPort_13[5:0]), //o
    .io_recoveryPort_14  (cpuClockingArea_aRAT_io_recoveryPort_14[5:0]), //o
    .io_recoveryPort_15  (cpuClockingArea_aRAT_io_recoveryPort_15[5:0]), //o
    .io_recoveryPort_16  (cpuClockingArea_aRAT_io_recoveryPort_16[5:0]), //o
    .io_recoveryPort_17  (cpuClockingArea_aRAT_io_recoveryPort_17[5:0]), //o
    .io_recoveryPort_18  (cpuClockingArea_aRAT_io_recoveryPort_18[5:0]), //o
    .io_recoveryPort_19  (cpuClockingArea_aRAT_io_recoveryPort_19[5:0]), //o
    .io_recoveryPort_20  (cpuClockingArea_aRAT_io_recoveryPort_20[5:0]), //o
    .io_recoveryPort_21  (cpuClockingArea_aRAT_io_recoveryPort_21[5:0]), //o
    .io_recoveryPort_22  (cpuClockingArea_aRAT_io_recoveryPort_22[5:0]), //o
    .io_recoveryPort_23  (cpuClockingArea_aRAT_io_recoveryPort_23[5:0]), //o
    .io_recoveryPort_24  (cpuClockingArea_aRAT_io_recoveryPort_24[5:0]), //o
    .io_recoveryPort_25  (cpuClockingArea_aRAT_io_recoveryPort_25[5:0]), //o
    .io_recoveryPort_26  (cpuClockingArea_aRAT_io_recoveryPort_26[5:0]), //o
    .io_recoveryPort_27  (cpuClockingArea_aRAT_io_recoveryPort_27[5:0]), //o
    .io_recoveryPort_28  (cpuClockingArea_aRAT_io_recoveryPort_28[5:0]), //o
    .io_recoveryPort_29  (cpuClockingArea_aRAT_io_recoveryPort_29[5:0]), //o
    .io_recoveryPort_30  (cpuClockingArea_aRAT_io_recoveryPort_30[5:0]), //o
    .io_recoveryPort_31  (cpuClockingArea_aRAT_io_recoveryPort_31[5:0]), //o
    .aclk                (aclk                                        ), //i
    .aresetn             (aresetn                                     )  //i
  );
  FreeList cpuClockingArea_freeList (
    .io_dispatch_disPatchNum (cpuClockingArea_areaFlushReset_dispatcher_io_freelist_disPatchNum[1:0]), //i
    .io_dispatch_availMask   (cpuClockingArea_freeList_io_dispatch_availMask[1:0]                   ), //o
    .io_dispatch_prfIdx_0    (cpuClockingArea_freeList_io_dispatch_prfIdx_0[5:0]                    ), //o
    .io_dispatch_prfIdx_1    (cpuClockingArea_freeList_io_dispatch_prfIdx_1[5:0]                    ), //o
    .io_retire_prfIdx_0      (cpuClockingArea_rob_io_retireFreeList_prfIdx_0[5:0]                   ), //i
    .io_retire_prfIdx_1      (cpuClockingArea_rob_io_retireFreeList_prfIdx_1[5:0]                   ), //i
    .io_retire_writeNum      (cpuClockingArea_rob_io_retireFreeList_writeNum[1:0]                   ), //i
    .io_retire_delayedFlush  (cpuClockingArea_rob_io_retireFreeList_delayedFlush                    ), //i
    .aclk                    (aclk                                                                  ), //i
    .aresetn                 (aresetn                                                               )  //i
  );
  PC cpuClockingArea_pc (
    .io_iCacheFeed_0_valid                            (cpuClockingArea_pc_io_iCacheFeed_0_valid                             ), //o
    .io_iCacheFeed_0_ready                            (cpuClockingArea_iCache_io_input_0_ready                              ), //i
    .io_iCacheFeed_0_payload_address                  (cpuClockingArea_pc_io_iCacheFeed_0_payload_address[31:0]             ), //o
    .io_iCacheFeed_0_payload_size                     (cpuClockingArea_pc_io_iCacheFeed_0_payload_size[3:0]                 ), //o
    .io_iCacheFeed_0_payload_branchInfo_predictPC     (cpuClockingArea_pc_io_iCacheFeed_0_payload_branchInfo_predictPC[31:0]), //o
    .io_iCacheFeed_0_payload_branchInfo_predictResult (cpuClockingArea_pc_io_iCacheFeed_0_payload_branchInfo_predictResult  ), //o
    .io_iCacheFeed_1_valid                            (cpuClockingArea_pc_io_iCacheFeed_1_valid                             ), //o
    .io_iCacheFeed_1_ready                            (cpuClockingArea_iCache_io_input_1_ready                              ), //i
    .io_iCacheFeed_1_payload_address                  (cpuClockingArea_pc_io_iCacheFeed_1_payload_address[31:0]             ), //o
    .io_iCacheFeed_1_payload_size                     (cpuClockingArea_pc_io_iCacheFeed_1_payload_size[3:0]                 ), //o
    .io_iCacheFeed_1_payload_branchInfo_predictPC     (cpuClockingArea_pc_io_iCacheFeed_1_payload_branchInfo_predictPC[31:0]), //o
    .io_iCacheFeed_1_payload_branchInfo_predictResult (cpuClockingArea_pc_io_iCacheFeed_1_payload_branchInfo_predictResult  ), //o
    .io_pc_0_valid                                    (cpuClockingArea_pc_io_pc_0_valid                                     ), //o
    .io_pc_0_payload                                  (cpuClockingArea_pc_io_pc_0_payload[31:0]                             ), //o
    .io_pc_1_valid                                    (cpuClockingArea_pc_io_pc_1_valid                                     ), //o
    .io_pc_1_payload                                  (cpuClockingArea_pc_io_pc_1_payload[31:0]                             ), //o
    .io_npc_0_valid                                   (cpuClockingArea_nextLinePredictor_io_npc_0_valid                     ), //i
    .io_npc_0_payload                                 (cpuClockingArea_nextLinePredictor_io_npc_0_payload[31:0]             ), //i
    .io_npc_1_valid                                   (cpuClockingArea_nextLinePredictor_io_npc_1_valid                     ), //i
    .io_npc_1_payload                                 (cpuClockingArea_nextLinePredictor_io_npc_1_payload[31:0]             ), //i
    .io_branchInfo_0_predictPC                        (cpuClockingArea_nextLinePredictor_io_branchInfo_0_predictPC[31:0]    ), //i
    .io_branchInfo_0_predictResult                    (cpuClockingArea_nextLinePredictor_io_branchInfo_0_predictResult      ), //i
    .io_branchInfo_1_predictPC                        (cpuClockingArea_nextLinePredictor_io_branchInfo_1_predictPC[31:0]    ), //i
    .io_branchInfo_1_predictResult                    (cpuClockingArea_nextLinePredictor_io_branchInfo_1_predictResult      ), //i
    .io_flush                                         (cpuClockingArea_rob_io_flush                                         ), //i
    .io_redirectPC                                    (cpuClockingArea_rob_io_redirectPC[31:0]                              ), //i
    .aclk                                             (aclk                                                                 ), //i
    .aresetn                                          (aresetn                                                              )  //i
  );
  NextLinePredictor cpuClockingArea_nextLinePredictor (
    .io_pc_0_valid                       (cpuClockingArea_pc_io_pc_0_valid                                 ), //i
    .io_pc_0_payload                     (cpuClockingArea_pc_io_pc_0_payload[31:0]                         ), //i
    .io_pc_1_valid                       (cpuClockingArea_pc_io_pc_1_valid                                 ), //i
    .io_pc_1_payload                     (cpuClockingArea_pc_io_pc_1_payload[31:0]                         ), //i
    .io_npc_0_valid                      (cpuClockingArea_nextLinePredictor_io_npc_0_valid                 ), //o
    .io_npc_0_payload                    (cpuClockingArea_nextLinePredictor_io_npc_0_payload[31:0]         ), //o
    .io_npc_1_valid                      (cpuClockingArea_nextLinePredictor_io_npc_1_valid                 ), //o
    .io_npc_1_payload                    (cpuClockingArea_nextLinePredictor_io_npc_1_payload[31:0]         ), //o
    .io_branchInfo_0_predictPC           (cpuClockingArea_nextLinePredictor_io_branchInfo_0_predictPC[31:0]), //o
    .io_branchInfo_0_predictResult       (cpuClockingArea_nextLinePredictor_io_branchInfo_0_predictResult  ), //o
    .io_branchInfo_1_predictPC           (cpuClockingArea_nextLinePredictor_io_branchInfo_1_predictPC[31:0]), //o
    .io_branchInfo_1_predictResult       (cpuClockingArea_nextLinePredictor_io_branchInfo_1_predictResult  ), //o
    .io_updateInfo_0_valid               (cpuClockingArea_rob_io_updateBPU_0_valid                         ), //i
    .io_updateInfo_0_payload_pc          (cpuClockingArea_rob_io_updateBPU_0_payload_pc[31:0]              ), //i
    .io_updateInfo_0_payload_isJumpInst  (cpuClockingArea_rob_io_updateBPU_0_payload_isJumpInst            ), //i
    .io_updateInfo_0_payload_taken       (cpuClockingArea_rob_io_updateBPU_0_payload_taken                 ), //i
    .io_updateInfo_0_payload_predictFail (cpuClockingArea_rob_io_updateBPU_0_payload_predictFail           ), //i
    .io_updateInfo_0_payload_target      (cpuClockingArea_rob_io_updateBPU_0_payload_target[31:0]          ), //i
    .io_updateInfo_1_valid               (cpuClockingArea_rob_io_updateBPU_1_valid                         ), //i
    .io_updateInfo_1_payload_pc          (cpuClockingArea_rob_io_updateBPU_1_payload_pc[31:0]              ), //i
    .io_updateInfo_1_payload_isJumpInst  (cpuClockingArea_rob_io_updateBPU_1_payload_isJumpInst            ), //i
    .io_updateInfo_1_payload_taken       (cpuClockingArea_rob_io_updateBPU_1_payload_taken                 ), //i
    .io_updateInfo_1_payload_predictFail (cpuClockingArea_rob_io_updateBPU_1_payload_predictFail           ), //i
    .io_updateInfo_1_payload_target      (cpuClockingArea_rob_io_updateBPU_1_payload_target[31:0]          )  //i
  );
  ICache cpuClockingArea_iCache (
    .io_input_0_valid                            (cpuClockingArea_pc_io_iCacheFeed_0_valid                             ), //i
    .io_input_0_ready                            (cpuClockingArea_iCache_io_input_0_ready                              ), //o
    .io_input_0_payload_address                  (cpuClockingArea_pc_io_iCacheFeed_0_payload_address[31:0]             ), //i
    .io_input_0_payload_size                     (cpuClockingArea_pc_io_iCacheFeed_0_payload_size[3:0]                 ), //i
    .io_input_0_payload_branchInfo_predictPC     (cpuClockingArea_pc_io_iCacheFeed_0_payload_branchInfo_predictPC[31:0]), //i
    .io_input_0_payload_branchInfo_predictResult (cpuClockingArea_pc_io_iCacheFeed_0_payload_branchInfo_predictResult  ), //i
    .io_input_1_valid                            (cpuClockingArea_pc_io_iCacheFeed_1_valid                             ), //i
    .io_input_1_ready                            (cpuClockingArea_iCache_io_input_1_ready                              ), //o
    .io_input_1_payload_address                  (cpuClockingArea_pc_io_iCacheFeed_1_payload_address[31:0]             ), //i
    .io_input_1_payload_size                     (cpuClockingArea_pc_io_iCacheFeed_1_payload_size[3:0]                 ), //i
    .io_input_1_payload_branchInfo_predictPC     (cpuClockingArea_pc_io_iCacheFeed_1_payload_branchInfo_predictPC[31:0]), //i
    .io_input_1_payload_branchInfo_predictResult (cpuClockingArea_pc_io_iCacheFeed_1_payload_branchInfo_predictResult  ), //i
    .io_output_allowMask                         (cpuClockingArea_areaFlushReset_instQueue_io_in_allowMask[1:0]        ), //i
    .io_output_availMask                         (cpuClockingArea_iCache_io_output_availMask[1:0]                      ), //o
    .io_output_info_0_inst                       (cpuClockingArea_iCache_io_output_info_0_inst[31:0]                   ), //o
    .io_output_info_0_branchInfo_predictPC       (cpuClockingArea_iCache_io_output_info_0_branchInfo_predictPC[31:0]   ), //o
    .io_output_info_0_branchInfo_predictResult   (cpuClockingArea_iCache_io_output_info_0_branchInfo_predictResult     ), //o
    .io_output_info_0_exceptionInfo_exception    (cpuClockingArea_iCache_io_output_info_0_exceptionInfo_exception      ), //o
    .io_output_info_0_exceptionInfo_eCode        (cpuClockingArea_iCache_io_output_info_0_exceptionInfo_eCode[5:0]     ), //o
    .io_output_info_0_exceptionInfo_eSubCode     (cpuClockingArea_iCache_io_output_info_0_exceptionInfo_eSubCode       ), //o
    .io_output_info_0_pc                         (cpuClockingArea_iCache_io_output_info_0_pc[31:0]                     ), //o
    .io_output_info_1_inst                       (cpuClockingArea_iCache_io_output_info_1_inst[31:0]                   ), //o
    .io_output_info_1_branchInfo_predictPC       (cpuClockingArea_iCache_io_output_info_1_branchInfo_predictPC[31:0]   ), //o
    .io_output_info_1_branchInfo_predictResult   (cpuClockingArea_iCache_io_output_info_1_branchInfo_predictResult     ), //o
    .io_output_info_1_exceptionInfo_exception    (cpuClockingArea_iCache_io_output_info_1_exceptionInfo_exception      ), //o
    .io_output_info_1_exceptionInfo_eCode        (cpuClockingArea_iCache_io_output_info_1_exceptionInfo_eCode[5:0]     ), //o
    .io_output_info_1_exceptionInfo_eSubCode     (cpuClockingArea_iCache_io_output_info_1_exceptionInfo_eSubCode       ), //o
    .io_output_info_1_pc                         (cpuClockingArea_iCache_io_output_info_1_pc[31:0]                     ), //o
    .io_tlb_hit                                  (cpuClockingArea_tlb_io_iCacheReq_hit                                 ), //i
    .io_tlb_pageInfo_ppn                         (cpuClockingArea_tlb_io_iCacheReq_pageInfo_ppn[19:0]                  ), //i
    .io_tlb_pageInfo_plv                         (cpuClockingArea_tlb_io_iCacheReq_pageInfo_plv[1:0]                   ), //i
    .io_tlb_pageInfo_mat                         (cpuClockingArea_tlb_io_iCacheReq_pageInfo_mat[1:0]                   ), //i
    .io_tlb_pageInfo_d                           (cpuClockingArea_tlb_io_iCacheReq_pageInfo_d                          ), //i
    .io_tlb_pageInfo_v                           (cpuClockingArea_tlb_io_iCacheReq_pageInfo_v                          ), //i
    .io_tlb_virtPageNumber                       (cpuClockingArea_iCache_io_tlb_virtPageNumber[19:0]                   ), //o
    ._zz_when_Cache_l83                          (cpuClockingArea_csr__zz_when_Cache_l83[1:0]                          ), //i
    .io_ctrl_busy                                (cpuClockingArea_iCache_io_ctrl_busy                                  ), //o
    .io_ctrl_stall                               (cpuClockingArea_memService_io_iCacheCtrl_stall                       ), //i
    .io_ctrl_cacopVA                             (cpuClockingArea_memService_io_iCacheCtrl_cacopVA[31:0]               ), //i
    .io_ctrl_cacopStoreTag                       (cpuClockingArea_memService_io_iCacheCtrl_cacopStoreTag               ), //i
    .io_ctrl_cacopIndexInvalidate                (cpuClockingArea_memService_io_iCacheCtrl_cacopIndexInvalidate        ), //i
    .io_ctrl_cacopHitInvalidate                  (cpuClockingArea_memService_io_iCacheCtrl_cacopHitInvalidate          ), //i
    .io_flush                                    (cpuClockingArea_rob_io_flush                                         ), //i
    .io_badv_vaddr                               (cpuClockingArea_iCache_io_badv_vaddr[31:0]                           ), //o
    .io_badv_wen                                 (cpuClockingArea_iCache_io_badv_wen                                   ), //o
    .io_axi_arid                                 (cpuClockingArea_iCache_io_axi_arid[3:0]                              ), //o
    .io_axi_araddr                               (cpuClockingArea_iCache_io_axi_araddr[31:0]                           ), //o
    .io_axi_arlen                                (cpuClockingArea_iCache_io_axi_arlen[7:0]                             ), //o
    .io_axi_arsize                               (cpuClockingArea_iCache_io_axi_arsize[2:0]                            ), //o
    .io_axi_arburst                              (cpuClockingArea_iCache_io_axi_arburst[1:0]                           ), //o
    .io_axi_arlock                               (cpuClockingArea_iCache_io_axi_arlock[1:0]                            ), //o
    .io_axi_arcache                              (cpuClockingArea_iCache_io_axi_arcache[3:0]                           ), //o
    .io_axi_arprot                               (cpuClockingArea_iCache_io_axi_arprot[2:0]                            ), //o
    .io_axi_arvalid                              (cpuClockingArea_iCache_io_axi_arvalid                                ), //o
    .io_axi_arready                              (cpuClockingArea_arbiter_io_iCache_arready                            ), //i
    .io_axi_rid                                  (cpuClockingArea_arbiter_io_iCache_rid[3:0]                           ), //i
    .io_axi_rdata                                (cpuClockingArea_arbiter_io_iCache_rdata[31:0]                        ), //i
    .io_axi_rresp                                (cpuClockingArea_arbiter_io_iCache_rresp[1:0]                         ), //i
    .io_axi_rlast                                (cpuClockingArea_arbiter_io_iCache_rlast                              ), //i
    .io_axi_rvalid                               (cpuClockingArea_arbiter_io_iCache_rvalid                             ), //i
    .io_axi_rready                               (cpuClockingArea_iCache_io_axi_rready                                 ), //o
    .aclk                                        (aclk                                                                 ), //i
    .aresetn                                     (aresetn                                                              )  //i
  );
  DCache cpuClockingArea_fuLSU (
    .io_input_valid                               (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_valid                              ), //i
    .io_input_ready                               (cpuClockingArea_fuLSU_io_input_ready                                                             ), //o
    .io_input_payload_src1                        (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_src1[31:0]                 ), //i
    .io_input_payload_src2                        (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_src2[31:0]                 ), //i
    .io_input_payload_src3                        (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_src3[31:0]                 ), //i
    .io_input_payload_robIdx                      (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_robIdx[4:0]                ), //i
    .io_input_payload_branchResult_targetPC       (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_branchResult_targetPC[31:0]), //i
    .io_input_payload_branchResult_branchResult   (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_branchResult_branchResult  ), //i
    .io_input_payload_branchResult_predictFail    (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_branchResult_predictFail   ), //i
    .io_input_payload_exceptionInfo_exception     (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_exceptionInfo_exception    ), //i
    .io_input_payload_exceptionInfo_eCode         (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_exceptionInfo_eCode[5:0]   ), //i
    .io_input_payload_exceptionInfo_eSubCode      (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode     ), //i
    .io_input_payload_pc                          (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_pc[31:0]                   ), //i
    .io_input_payload_prd                         (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_prd[5:0]                   ), //i
    .io_input_payload_uop_lsuOp                   (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp[3:0]             ), //i
    .io_input_payload_uop_lsuCoOp                 (toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuCoOp[4:0]           ), //i
    .io_output_valid                              (cpuClockingArea_fuLSU_io_output_valid                                                            ), //o
    .io_output_ready                              (cpuClockingArea_fuLSU_io_output_ready                                                            ), //i
    .io_output_payload_robIdx                     (cpuClockingArea_fuLSU_io_output_payload_robIdx[4:0]                                              ), //o
    .io_output_payload_data                       (cpuClockingArea_fuLSU_io_output_payload_data[31:0]                                               ), //o
    .io_output_payload_prd                        (cpuClockingArea_fuLSU_io_output_payload_prd[5:0]                                                 ), //o
    .io_output_payload_branchResult_targetPC      (cpuClockingArea_fuLSU_io_output_payload_branchResult_targetPC[31:0]                              ), //o
    .io_output_payload_branchResult_branchResult  (cpuClockingArea_fuLSU_io_output_payload_branchResult_branchResult                                ), //o
    .io_output_payload_branchResult_predictFail   (cpuClockingArea_fuLSU_io_output_payload_branchResult_predictFail                                 ), //o
    .io_output_payload_exceptionInfo_exception    (cpuClockingArea_fuLSU_io_output_payload_exceptionInfo_exception                                  ), //o
    .io_output_payload_exceptionInfo_eCode        (cpuClockingArea_fuLSU_io_output_payload_exceptionInfo_eCode[5:0]                                 ), //o
    .io_output_payload_exceptionInfo_eSubCode     (cpuClockingArea_fuLSU_io_output_payload_exceptionInfo_eSubCode                                   ), //o
    .io_wakeOut_0_valid                           (cpuClockingArea_fuLSU_io_wakeOut_0_valid                                                         ), //o
    .io_wakeOut_0_payload                         (cpuClockingArea_fuLSU_io_wakeOut_0_payload[5:0]                                                  ), //o
    .io_wakeOut_1_valid                           (cpuClockingArea_fuLSU_io_wakeOut_1_valid                                                         ), //o
    .io_wakeOut_1_payload                         (cpuClockingArea_fuLSU_io_wakeOut_1_payload[5:0]                                                  ), //o
    .io_retireComm_robIdx_0                       (cpuClockingArea_rob_io_retireLSU_robIdx_0[4:0]                                                   ), //i
    .io_retireComm_robIdx_1                       (cpuClockingArea_rob_io_retireLSU_robIdx_1[4:0]                                                   ), //i
    .io_retireComm_allowRetire_0                  (cpuClockingArea_rob_io_retireLSU_allowRetire_0                                                   ), //i
    .io_retireComm_allowRetire_1                  (cpuClockingArea_rob_io_retireLSU_allowRetire_1                                                   ), //i
    .io_tlb_hit                                   (cpuClockingArea_tlb_io_dCacheReq_hit                                                             ), //i
    .io_tlb_pageInfo_ppn                          (cpuClockingArea_tlb_io_dCacheReq_pageInfo_ppn[19:0]                                              ), //i
    .io_tlb_pageInfo_plv                          (cpuClockingArea_tlb_io_dCacheReq_pageInfo_plv[1:0]                                               ), //i
    .io_tlb_pageInfo_mat                          (cpuClockingArea_tlb_io_dCacheReq_pageInfo_mat[1:0]                                               ), //i
    .io_tlb_pageInfo_d                            (cpuClockingArea_tlb_io_dCacheReq_pageInfo_d                                                      ), //i
    .io_tlb_pageInfo_v                            (cpuClockingArea_tlb_io_dCacheReq_pageInfo_v                                                      ), //i
    .io_tlb_virtPageNumber                        (cpuClockingArea_fuLSU_io_tlb_virtPageNumber[19:0]                                                ), //o
    ._zz_when_LSU_l217                            (cpuClockingArea_csr__zz_when_Cache_l83[1:0]                                                      ), //i
    .io_llBitComm_actualAddr                      (cpuClockingArea_csr_io_llBitComm_actualAddr[31:0]                                                ), //i
    .io_llBitComm_toUpdateAddr                    (cpuClockingArea_fuLSU_io_llBitComm_toUpdateAddr[31:0]                                            ), //o
    .io_llBitComm_wen                             (cpuClockingArea_fuLSU_io_llBitComm_wen                                                           ), //o
    ._zz_scMatchHit                               (cpuClockingArea_csr__zz_scMatchHit                                                               ), //i
    .io_ctrl_busy                                 (cpuClockingArea_fuLSU_io_ctrl_busy                                                               ), //o
    .io_ctrl_stall                                (cpuClockingArea_memService_io_dCacheCtrl_stall                                                   ), //i
    .io_ctrl_cacopVA                              (cpuClockingArea_memService_io_dCacheCtrl_cacopVA[31:0]                                           ), //i
    .io_ctrl_cacopStoreTag                        (cpuClockingArea_memService_io_dCacheCtrl_cacopStoreTag                                           ), //i
    .io_ctrl_cacopIndexInvalidate                 (cpuClockingArea_memService_io_dCacheCtrl_cacopIndexInvalidate                                    ), //i
    .io_ctrl_cacopHitInvalidate                   (cpuClockingArea_memService_io_dCacheCtrl_cacopHitInvalidate                                      ), //i
    .io_specialOpBufferUpdate_valid               (cpuClockingArea_fuLSU_io_specialOpBufferUpdate_valid                                             ), //o
    .io_specialOpBufferUpdate_payload_uop_lsuOp   (cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_uop_lsuOp[3:0]                            ), //o
    .io_specialOpBufferUpdate_payload_uop_lsuCoOp (cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_uop_lsuCoOp[4:0]                          ), //o
    .io_specialOpBufferUpdate_payload_vaddr       (cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_vaddr[31:0]                               ), //o
    .io_specialOpBufferUpdate_payload_asid        (cpuClockingArea_fuLSU_io_specialOpBufferUpdate_payload_asid[9:0]                                 ), //o
    .io_flush                                     (cpuClockingArea_rob_io_flush                                                                     ), //i
    .io_badv_robIdx                               (cpuClockingArea_fuLSU_io_badv_robIdx[4:0]                                                        ), //o
    .io_badv_vaddr                                (cpuClockingArea_fuLSU_io_badv_vaddr[31:0]                                                        ), //o
    .io_badv_wen                                  (cpuClockingArea_fuLSU_io_badv_wen                                                                ), //o
    .io_axi_arid                                  (cpuClockingArea_fuLSU_io_axi_arid[3:0]                                                           ), //o
    .io_axi_araddr                                (cpuClockingArea_fuLSU_io_axi_araddr[31:0]                                                        ), //o
    .io_axi_arlen                                 (cpuClockingArea_fuLSU_io_axi_arlen[7:0]                                                          ), //o
    .io_axi_arsize                                (cpuClockingArea_fuLSU_io_axi_arsize[2:0]                                                         ), //o
    .io_axi_arburst                               (cpuClockingArea_fuLSU_io_axi_arburst[1:0]                                                        ), //o
    .io_axi_arlock                                (cpuClockingArea_fuLSU_io_axi_arlock[1:0]                                                         ), //o
    .io_axi_arcache                               (cpuClockingArea_fuLSU_io_axi_arcache[3:0]                                                        ), //o
    .io_axi_arprot                                (cpuClockingArea_fuLSU_io_axi_arprot[2:0]                                                         ), //o
    .io_axi_arvalid                               (cpuClockingArea_fuLSU_io_axi_arvalid                                                             ), //o
    .io_axi_arready                               (cpuClockingArea_arbiter_io_dCache_arready                                                        ), //i
    .io_axi_rid                                   (cpuClockingArea_arbiter_io_dCache_rid[3:0]                                                       ), //i
    .io_axi_rdata                                 (cpuClockingArea_arbiter_io_dCache_rdata[31:0]                                                    ), //i
    .io_axi_rresp                                 (cpuClockingArea_arbiter_io_dCache_rresp[1:0]                                                     ), //i
    .io_axi_rlast                                 (cpuClockingArea_arbiter_io_dCache_rlast                                                          ), //i
    .io_axi_rvalid                                (cpuClockingArea_arbiter_io_dCache_rvalid                                                         ), //i
    .io_axi_rready                                (cpuClockingArea_fuLSU_io_axi_rready                                                              ), //o
    .io_axi_awid                                  (cpuClockingArea_fuLSU_io_axi_awid[3:0]                                                           ), //o
    .io_axi_awaddr                                (cpuClockingArea_fuLSU_io_axi_awaddr[31:0]                                                        ), //o
    .io_axi_awlen                                 (cpuClockingArea_fuLSU_io_axi_awlen[7:0]                                                          ), //o
    .io_axi_awsize                                (cpuClockingArea_fuLSU_io_axi_awsize[2:0]                                                         ), //o
    .io_axi_awburst                               (cpuClockingArea_fuLSU_io_axi_awburst[1:0]                                                        ), //o
    .io_axi_awlock                                (cpuClockingArea_fuLSU_io_axi_awlock[1:0]                                                         ), //o
    .io_axi_awcache                               (cpuClockingArea_fuLSU_io_axi_awcache[3:0]                                                        ), //o
    .io_axi_awprot                                (cpuClockingArea_fuLSU_io_axi_awprot[2:0]                                                         ), //o
    .io_axi_awvalid                               (cpuClockingArea_fuLSU_io_axi_awvalid                                                             ), //o
    .io_axi_awready                               (cpuClockingArea_arbiter_io_dCache_awready                                                        ), //i
    .io_axi_wid                                   (cpuClockingArea_fuLSU_io_axi_wid[3:0]                                                            ), //o
    .io_axi_wdata                                 (cpuClockingArea_fuLSU_io_axi_wdata[31:0]                                                         ), //o
    .io_axi_wstrb                                 (cpuClockingArea_fuLSU_io_axi_wstrb[3:0]                                                          ), //o
    .io_axi_wlast                                 (cpuClockingArea_fuLSU_io_axi_wlast                                                               ), //o
    .io_axi_wvalid                                (cpuClockingArea_fuLSU_io_axi_wvalid                                                              ), //o
    .io_axi_wready                                (cpuClockingArea_arbiter_io_dCache_wready                                                         ), //i
    .io_axi_bid                                   (cpuClockingArea_arbiter_io_dCache_bid[3:0]                                                       ), //i
    .io_axi_bresp                                 (cpuClockingArea_arbiter_io_dCache_bresp[1:0]                                                     ), //i
    .io_axi_bvalid                                (cpuClockingArea_arbiter_io_dCache_bvalid                                                         ), //i
    .io_axi_bready                                (cpuClockingArea_fuLSU_io_axi_bready                                                              ), //o
    .io_storeData                                 (cpuClockingArea_fuLSU_io_storeData[31:0]                                                         ), //o
    .io_storeMask                                 (cpuClockingArea_fuLSU_io_storeMask[3:0]                                                          ), //o
    .io_loadMask                                  (cpuClockingArea_fuLSU_io_loadMask[3:0]                                                           ), //o
    .io_VAddr                                     (cpuClockingArea_fuLSU_io_VAddr[31:0]                                                             ), //o
    .io_PAddr                                     (cpuClockingArea_fuLSU_io_PAddr[31:0]                                                             ), //o
    .aclk                                         (aclk                                                                                             ), //i
    .aresetn                                      (aresetn                                                                                          )  //i
  );
  PRF cpuClockingArea_prf (
    .io_read_0_0_idx  (cpuClockingArea_areaFlushReset_roALU0_io_prf_0_idx[5:0]    ), //i
    .io_read_0_0_data (cpuClockingArea_prf_io_read_0_0_data[31:0]                 ), //o
    .io_read_0_1_idx  (cpuClockingArea_areaFlushReset_roALU0_io_prf_1_idx[5:0]    ), //i
    .io_read_0_1_data (cpuClockingArea_prf_io_read_0_1_data[31:0]                 ), //o
    .io_read_1_0_idx  (cpuClockingArea_areaFlushReset_roALU1_io_prf_0_idx[5:0]    ), //i
    .io_read_1_0_data (cpuClockingArea_prf_io_read_1_0_data[31:0]                 ), //o
    .io_read_1_1_idx  (cpuClockingArea_areaFlushReset_roALU1_io_prf_1_idx[5:0]    ), //i
    .io_read_1_1_data (cpuClockingArea_prf_io_read_1_1_data[31:0]                 ), //o
    .io_read_2_0_idx  (cpuClockingArea_areaFlushReset_roMULU_io_prf_0_idx[5:0]    ), //i
    .io_read_2_0_data (cpuClockingArea_prf_io_read_2_0_data[31:0]                 ), //o
    .io_read_2_1_idx  (cpuClockingArea_areaFlushReset_roMULU_io_prf_1_idx[5:0]    ), //i
    .io_read_2_1_data (cpuClockingArea_prf_io_read_2_1_data[31:0]                 ), //o
    .io_read_3_0_idx  (cpuClockingArea_areaFlushReset_roDIVU_io_prf_0_idx[5:0]    ), //i
    .io_read_3_0_data (cpuClockingArea_prf_io_read_3_0_data[31:0]                 ), //o
    .io_read_3_1_idx  (cpuClockingArea_areaFlushReset_roDIVU_io_prf_1_idx[5:0]    ), //i
    .io_read_3_1_data (cpuClockingArea_prf_io_read_3_1_data[31:0]                 ), //o
    .io_read_4_0_idx  (cpuClockingArea_areaFlushReset_roLSU_io_prf_0_idx[5:0]     ), //i
    .io_read_4_0_data (cpuClockingArea_prf_io_read_4_0_data[31:0]                 ), //o
    .io_read_4_1_idx  (cpuClockingArea_areaFlushReset_roLSU_io_prf_1_idx[5:0]     ), //i
    .io_read_4_1_data (cpuClockingArea_prf_io_read_4_1_data[31:0]                 ), //o
    .io_write_0_idx   (cpuClockingArea_areaFlushReset_commitALU0_io_prf_idx[5:0]  ), //i
    .io_write_0_data  (cpuClockingArea_areaFlushReset_commitALU0_io_prf_data[31:0]), //i
    .io_write_1_idx   (cpuClockingArea_areaFlushReset_commitALU1_io_prf_idx[5:0]  ), //i
    .io_write_1_data  (cpuClockingArea_areaFlushReset_commitALU1_io_prf_data[31:0]), //i
    .io_write_2_idx   (cpuClockingArea_areaFlushReset_commitMULU_io_prf_idx[5:0]  ), //i
    .io_write_2_data  (cpuClockingArea_areaFlushReset_commitMULU_io_prf_data[31:0]), //i
    .io_write_3_idx   (cpuClockingArea_areaFlushReset_commitDIVU_io_prf_idx[5:0]  ), //i
    .io_write_3_data  (cpuClockingArea_areaFlushReset_commitDIVU_io_prf_data[31:0]), //i
    .io_write_4_idx   (cpuClockingArea_areaFlushReset_commitLSU_io_prf_idx[5:0]   ), //i
    .io_write_4_data  (cpuClockingArea_areaFlushReset_commitLSU_io_prf_data[31:0] ), //i
    .io_debugRegs_0   (cpuClockingArea_prf_io_debugRegs_0[31:0]                   ), //o
    .io_debugRegs_1   (cpuClockingArea_prf_io_debugRegs_1[31:0]                   ), //o
    .io_debugRegs_2   (cpuClockingArea_prf_io_debugRegs_2[31:0]                   ), //o
    .io_debugRegs_3   (cpuClockingArea_prf_io_debugRegs_3[31:0]                   ), //o
    .io_debugRegs_4   (cpuClockingArea_prf_io_debugRegs_4[31:0]                   ), //o
    .io_debugRegs_5   (cpuClockingArea_prf_io_debugRegs_5[31:0]                   ), //o
    .io_debugRegs_6   (cpuClockingArea_prf_io_debugRegs_6[31:0]                   ), //o
    .io_debugRegs_7   (cpuClockingArea_prf_io_debugRegs_7[31:0]                   ), //o
    .io_debugRegs_8   (cpuClockingArea_prf_io_debugRegs_8[31:0]                   ), //o
    .io_debugRegs_9   (cpuClockingArea_prf_io_debugRegs_9[31:0]                   ), //o
    .io_debugRegs_10  (cpuClockingArea_prf_io_debugRegs_10[31:0]                  ), //o
    .io_debugRegs_11  (cpuClockingArea_prf_io_debugRegs_11[31:0]                  ), //o
    .io_debugRegs_12  (cpuClockingArea_prf_io_debugRegs_12[31:0]                  ), //o
    .io_debugRegs_13  (cpuClockingArea_prf_io_debugRegs_13[31:0]                  ), //o
    .io_debugRegs_14  (cpuClockingArea_prf_io_debugRegs_14[31:0]                  ), //o
    .io_debugRegs_15  (cpuClockingArea_prf_io_debugRegs_15[31:0]                  ), //o
    .io_debugRegs_16  (cpuClockingArea_prf_io_debugRegs_16[31:0]                  ), //o
    .io_debugRegs_17  (cpuClockingArea_prf_io_debugRegs_17[31:0]                  ), //o
    .io_debugRegs_18  (cpuClockingArea_prf_io_debugRegs_18[31:0]                  ), //o
    .io_debugRegs_19  (cpuClockingArea_prf_io_debugRegs_19[31:0]                  ), //o
    .io_debugRegs_20  (cpuClockingArea_prf_io_debugRegs_20[31:0]                  ), //o
    .io_debugRegs_21  (cpuClockingArea_prf_io_debugRegs_21[31:0]                  ), //o
    .io_debugRegs_22  (cpuClockingArea_prf_io_debugRegs_22[31:0]                  ), //o
    .io_debugRegs_23  (cpuClockingArea_prf_io_debugRegs_23[31:0]                  ), //o
    .io_debugRegs_24  (cpuClockingArea_prf_io_debugRegs_24[31:0]                  ), //o
    .io_debugRegs_25  (cpuClockingArea_prf_io_debugRegs_25[31:0]                  ), //o
    .io_debugRegs_26  (cpuClockingArea_prf_io_debugRegs_26[31:0]                  ), //o
    .io_debugRegs_27  (cpuClockingArea_prf_io_debugRegs_27[31:0]                  ), //o
    .io_debugRegs_28  (cpuClockingArea_prf_io_debugRegs_28[31:0]                  ), //o
    .io_debugRegs_29  (cpuClockingArea_prf_io_debugRegs_29[31:0]                  ), //o
    .io_debugRegs_30  (cpuClockingArea_prf_io_debugRegs_30[31:0]                  ), //o
    .io_debugRegs_31  (cpuClockingArea_prf_io_debugRegs_31[31:0]                  ), //o
    .io_debugRegs_32  (cpuClockingArea_prf_io_debugRegs_32[31:0]                  ), //o
    .io_debugRegs_33  (cpuClockingArea_prf_io_debugRegs_33[31:0]                  ), //o
    .io_debugRegs_34  (cpuClockingArea_prf_io_debugRegs_34[31:0]                  ), //o
    .io_debugRegs_35  (cpuClockingArea_prf_io_debugRegs_35[31:0]                  ), //o
    .io_debugRegs_36  (cpuClockingArea_prf_io_debugRegs_36[31:0]                  ), //o
    .io_debugRegs_37  (cpuClockingArea_prf_io_debugRegs_37[31:0]                  ), //o
    .io_debugRegs_38  (cpuClockingArea_prf_io_debugRegs_38[31:0]                  ), //o
    .io_debugRegs_39  (cpuClockingArea_prf_io_debugRegs_39[31:0]                  ), //o
    .io_debugRegs_40  (cpuClockingArea_prf_io_debugRegs_40[31:0]                  ), //o
    .io_debugRegs_41  (cpuClockingArea_prf_io_debugRegs_41[31:0]                  ), //o
    .io_debugRegs_42  (cpuClockingArea_prf_io_debugRegs_42[31:0]                  ), //o
    .io_debugRegs_43  (cpuClockingArea_prf_io_debugRegs_43[31:0]                  ), //o
    .io_debugRegs_44  (cpuClockingArea_prf_io_debugRegs_44[31:0]                  ), //o
    .io_debugRegs_45  (cpuClockingArea_prf_io_debugRegs_45[31:0]                  ), //o
    .io_debugRegs_46  (cpuClockingArea_prf_io_debugRegs_46[31:0]                  ), //o
    .io_debugRegs_47  (cpuClockingArea_prf_io_debugRegs_47[31:0]                  ), //o
    .io_debugRegs_48  (cpuClockingArea_prf_io_debugRegs_48[31:0]                  ), //o
    .io_debugRegs_49  (cpuClockingArea_prf_io_debugRegs_49[31:0]                  ), //o
    .io_debugRegs_50  (cpuClockingArea_prf_io_debugRegs_50[31:0]                  ), //o
    .io_debugRegs_51  (cpuClockingArea_prf_io_debugRegs_51[31:0]                  ), //o
    .io_debugRegs_52  (cpuClockingArea_prf_io_debugRegs_52[31:0]                  ), //o
    .io_debugRegs_53  (cpuClockingArea_prf_io_debugRegs_53[31:0]                  ), //o
    .io_debugRegs_54  (cpuClockingArea_prf_io_debugRegs_54[31:0]                  ), //o
    .io_debugRegs_55  (cpuClockingArea_prf_io_debugRegs_55[31:0]                  ), //o
    .io_debugRegs_56  (cpuClockingArea_prf_io_debugRegs_56[31:0]                  ), //o
    .io_debugRegs_57  (cpuClockingArea_prf_io_debugRegs_57[31:0]                  ), //o
    .io_debugRegs_58  (cpuClockingArea_prf_io_debugRegs_58[31:0]                  ), //o
    .io_debugRegs_59  (cpuClockingArea_prf_io_debugRegs_59[31:0]                  ), //o
    .io_debugRegs_60  (cpuClockingArea_prf_io_debugRegs_60[31:0]                  ), //o
    .io_debugRegs_61  (cpuClockingArea_prf_io_debugRegs_61[31:0]                  ), //o
    .io_debugRegs_62  (cpuClockingArea_prf_io_debugRegs_62[31:0]                  ), //o
    .io_debugRegs_63  (cpuClockingArea_prf_io_debugRegs_63[31:0]                  ), //o
    .aclk             (aclk                                                       ), //i
    .aresetn          (aresetn                                                    )  //i
  );
  ROB cpuClockingArea_rob (
    .io_dispatch_allowMask                           (cpuClockingArea_areaFlushReset_dispatcher_io_rob_allowMask[1:0]             ), //i
    .io_dispatch_availMask                           (cpuClockingArea_rob_io_dispatch_availMask[1:0]                              ), //o
    .io_dispatch_robIdx_0                            (cpuClockingArea_rob_io_dispatch_robIdx_0[4:0]                               ), //o
    .io_dispatch_robIdx_1                            (cpuClockingArea_rob_io_dispatch_robIdx_1[4:0]                               ), //o
    .io_dispatch_pc_0                                (cpuClockingArea_areaFlushReset_dispatcher_io_rob_pc_0[31:0]                 ), //i
    .io_dispatch_pc_1                                (cpuClockingArea_areaFlushReset_dispatcher_io_rob_pc_1[31:0]                 ), //i
    .io_dispatch_ard_0                               (cpuClockingArea_areaFlushReset_dispatcher_io_rob_ard_0[4:0]                 ), //i
    .io_dispatch_ard_1                               (cpuClockingArea_areaFlushReset_dispatcher_io_rob_ard_1[4:0]                 ), //i
    .io_dispatch_prd_0                               (cpuClockingArea_areaFlushReset_dispatcher_io_rob_prd_0[5:0]                 ), //i
    .io_dispatch_prd_1                               (cpuClockingArea_areaFlushReset_dispatcher_io_rob_prd_1[5:0]                 ), //i
    .io_dispatch_pprd_0                              (cpuClockingArea_areaFlushReset_dispatcher_io_rob_pprd_0[5:0]                ), //i
    .io_dispatch_pprd_1                              (cpuClockingArea_areaFlushReset_dispatcher_io_rob_pprd_1[5:0]                ), //i
    .io_dispatch_specialOp_0                         (cpuClockingArea_areaFlushReset_dispatcher_io_rob_specialOp_0[3:0]           ), //i
    .io_dispatch_specialOp_1                         (cpuClockingArea_areaFlushReset_dispatcher_io_rob_specialOp_1[3:0]           ), //i
    .io_commit_0_robIdx                              (cpuClockingArea_areaFlushReset_commitALU0_io_rob_robIdx[4:0]                ), //i
    .io_commit_0_branchResult_targetPC               (cpuClockingArea_areaFlushReset_commitALU0_io_rob_branchResult_targetPC[31:0]), //i
    .io_commit_0_branchResult_branchResult           (cpuClockingArea_areaFlushReset_commitALU0_io_rob_branchResult_branchResult  ), //i
    .io_commit_0_branchResult_predictFail            (cpuClockingArea_areaFlushReset_commitALU0_io_rob_branchResult_predictFail   ), //i
    .io_commit_0_exceptionInfo_exception             (cpuClockingArea_areaFlushReset_commitALU0_io_rob_exceptionInfo_exception    ), //i
    .io_commit_0_exceptionInfo_eCode                 (cpuClockingArea_areaFlushReset_commitALU0_io_rob_exceptionInfo_eCode[5:0]   ), //i
    .io_commit_0_exceptionInfo_eSubCode              (cpuClockingArea_areaFlushReset_commitALU0_io_rob_exceptionInfo_eSubCode     ), //i
    .io_commit_0_valid                               (cpuClockingArea_areaFlushReset_commitALU0_io_rob_valid                      ), //i
    .io_commit_1_robIdx                              (cpuClockingArea_areaFlushReset_commitALU1_io_rob_robIdx[4:0]                ), //i
    .io_commit_1_branchResult_targetPC               (cpuClockingArea_areaFlushReset_commitALU1_io_rob_branchResult_targetPC[31:0]), //i
    .io_commit_1_branchResult_branchResult           (cpuClockingArea_areaFlushReset_commitALU1_io_rob_branchResult_branchResult  ), //i
    .io_commit_1_branchResult_predictFail            (cpuClockingArea_areaFlushReset_commitALU1_io_rob_branchResult_predictFail   ), //i
    .io_commit_1_exceptionInfo_exception             (cpuClockingArea_areaFlushReset_commitALU1_io_rob_exceptionInfo_exception    ), //i
    .io_commit_1_exceptionInfo_eCode                 (cpuClockingArea_areaFlushReset_commitALU1_io_rob_exceptionInfo_eCode[5:0]   ), //i
    .io_commit_1_exceptionInfo_eSubCode              (cpuClockingArea_areaFlushReset_commitALU1_io_rob_exceptionInfo_eSubCode     ), //i
    .io_commit_1_valid                               (cpuClockingArea_areaFlushReset_commitALU1_io_rob_valid                      ), //i
    .io_commit_2_robIdx                              (cpuClockingArea_areaFlushReset_commitMULU_io_rob_robIdx[4:0]                ), //i
    .io_commit_2_branchResult_targetPC               (cpuClockingArea_areaFlushReset_commitMULU_io_rob_branchResult_targetPC[31:0]), //i
    .io_commit_2_branchResult_branchResult           (cpuClockingArea_areaFlushReset_commitMULU_io_rob_branchResult_branchResult  ), //i
    .io_commit_2_branchResult_predictFail            (cpuClockingArea_areaFlushReset_commitMULU_io_rob_branchResult_predictFail   ), //i
    .io_commit_2_exceptionInfo_exception             (cpuClockingArea_areaFlushReset_commitMULU_io_rob_exceptionInfo_exception    ), //i
    .io_commit_2_exceptionInfo_eCode                 (cpuClockingArea_areaFlushReset_commitMULU_io_rob_exceptionInfo_eCode[5:0]   ), //i
    .io_commit_2_exceptionInfo_eSubCode              (cpuClockingArea_areaFlushReset_commitMULU_io_rob_exceptionInfo_eSubCode     ), //i
    .io_commit_2_valid                               (cpuClockingArea_areaFlushReset_commitMULU_io_rob_valid                      ), //i
    .io_commit_3_robIdx                              (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_robIdx[4:0]                ), //i
    .io_commit_3_branchResult_targetPC               (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_branchResult_targetPC[31:0]), //i
    .io_commit_3_branchResult_branchResult           (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_branchResult_branchResult  ), //i
    .io_commit_3_branchResult_predictFail            (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_branchResult_predictFail   ), //i
    .io_commit_3_exceptionInfo_exception             (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_exceptionInfo_exception    ), //i
    .io_commit_3_exceptionInfo_eCode                 (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_exceptionInfo_eCode[5:0]   ), //i
    .io_commit_3_exceptionInfo_eSubCode              (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_exceptionInfo_eSubCode     ), //i
    .io_commit_3_valid                               (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_valid                      ), //i
    .io_commit_4_robIdx                              (cpuClockingArea_areaFlushReset_commitLSU_io_rob_robIdx[4:0]                 ), //i
    .io_commit_4_branchResult_targetPC               (cpuClockingArea_areaFlushReset_commitLSU_io_rob_branchResult_targetPC[31:0] ), //i
    .io_commit_4_branchResult_branchResult           (cpuClockingArea_areaFlushReset_commitLSU_io_rob_branchResult_branchResult   ), //i
    .io_commit_4_branchResult_predictFail            (cpuClockingArea_areaFlushReset_commitLSU_io_rob_branchResult_predictFail    ), //i
    .io_commit_4_exceptionInfo_exception             (cpuClockingArea_areaFlushReset_commitLSU_io_rob_exceptionInfo_exception     ), //i
    .io_commit_4_exceptionInfo_eCode                 (cpuClockingArea_areaFlushReset_commitLSU_io_rob_exceptionInfo_eCode[5:0]    ), //i
    .io_commit_4_exceptionInfo_eSubCode              (cpuClockingArea_areaFlushReset_commitLSU_io_rob_exceptionInfo_eSubCode      ), //i
    .io_commit_4_valid                               (cpuClockingArea_areaFlushReset_commitLSU_io_rob_valid                       ), //i
    .io_retireARAT_0_ard                             (cpuClockingArea_rob_io_retireARAT_0_ard[4:0]                                ), //o
    .io_retireARAT_0_prd                             (cpuClockingArea_rob_io_retireARAT_0_prd[5:0]                                ), //o
    .io_retireARAT_0_wen                             (cpuClockingArea_rob_io_retireARAT_0_wen                                     ), //o
    .io_retireARAT_1_ard                             (cpuClockingArea_rob_io_retireARAT_1_ard[4:0]                                ), //o
    .io_retireARAT_1_prd                             (cpuClockingArea_rob_io_retireARAT_1_prd[5:0]                                ), //o
    .io_retireARAT_1_wen                             (cpuClockingArea_rob_io_retireARAT_1_wen                                     ), //o
    .io_retireFreeList_prfIdx_0                      (cpuClockingArea_rob_io_retireFreeList_prfIdx_0[5:0]                         ), //o
    .io_retireFreeList_prfIdx_1                      (cpuClockingArea_rob_io_retireFreeList_prfIdx_1[5:0]                         ), //o
    .io_retireFreeList_writeNum                      (cpuClockingArea_rob_io_retireFreeList_writeNum[1:0]                         ), //o
    .io_retireFreeList_delayedFlush                  (cpuClockingArea_rob_io_retireFreeList_delayedFlush                          ), //o
    .io_retireLSU_robIdx_0                           (cpuClockingArea_rob_io_retireLSU_robIdx_0[4:0]                              ), //o
    .io_retireLSU_robIdx_1                           (cpuClockingArea_rob_io_retireLSU_robIdx_1[4:0]                              ), //o
    .io_retireLSU_allowRetire_0                      (cpuClockingArea_rob_io_retireLSU_allowRetire_0                              ), //o
    .io_retireLSU_allowRetire_1                      (cpuClockingArea_rob_io_retireLSU_allowRetire_1                              ), //o
    .io_wakeupMem                                    (cpuClockingArea_rob_io_wakeupMem                                            ), //o
    .io_updateBPU_0_valid                            (cpuClockingArea_rob_io_updateBPU_0_valid                                    ), //o
    .io_updateBPU_0_payload_pc                       (cpuClockingArea_rob_io_updateBPU_0_payload_pc[31:0]                         ), //o
    .io_updateBPU_0_payload_isJumpInst               (cpuClockingArea_rob_io_updateBPU_0_payload_isJumpInst                       ), //o
    .io_updateBPU_0_payload_taken                    (cpuClockingArea_rob_io_updateBPU_0_payload_taken                            ), //o
    .io_updateBPU_0_payload_predictFail              (cpuClockingArea_rob_io_updateBPU_0_payload_predictFail                      ), //o
    .io_updateBPU_0_payload_target                   (cpuClockingArea_rob_io_updateBPU_0_payload_target[31:0]                     ), //o
    .io_updateBPU_1_valid                            (cpuClockingArea_rob_io_updateBPU_1_valid                                    ), //o
    .io_updateBPU_1_payload_pc                       (cpuClockingArea_rob_io_updateBPU_1_payload_pc[31:0]                         ), //o
    .io_updateBPU_1_payload_isJumpInst               (cpuClockingArea_rob_io_updateBPU_1_payload_isJumpInst                       ), //o
    .io_updateBPU_1_payload_taken                    (cpuClockingArea_rob_io_updateBPU_1_payload_taken                            ), //o
    .io_updateBPU_1_payload_predictFail              (cpuClockingArea_rob_io_updateBPU_1_payload_predictFail                      ), //o
    .io_updateBPU_1_payload_target                   (cpuClockingArea_rob_io_updateBPU_1_payload_target[31:0]                     ), //o
    .io_csrCtrl_llBitUpdate                          (cpuClockingArea_rob_io_csrCtrl_llBitUpdate                                  ), //o
    .io_csrCtrl_writeCSR                             (cpuClockingArea_rob_io_csrCtrl_writeCSR                                     ), //o
    .io_csrCtrl_ertn                                 (cpuClockingArea_rob_io_csrCtrl_ertn                                         ), //o
    .io_csrCtrl_normalException                      (cpuClockingArea_rob_io_csrCtrl_normalException                              ), //o
    .io_csrCtrl_tlbrException                        (cpuClockingArea_rob_io_csrCtrl_tlbrException                                ), //o
    .io_csrCtrl_epc                                  (cpuClockingArea_rob_io_csrCtrl_epc[31:0]                                    ), //o
    .io_csrCtrl_eROBIdx                              (cpuClockingArea_rob_io_csrCtrl_eROBIdx[4:0]                                 ), //o
    .io_csrCtrl_eCode                                (cpuClockingArea_rob_io_csrCtrl_eCode[5:0]                                   ), //o
    .io_csrCtrl_eSubCode                             (cpuClockingArea_rob_io_csrCtrl_eSubCode                                     ), //o
    .io_csrCtrl_era                                  (cpuClockingArea_csr_io_ctrl_era[31:0]                                       ), //i
    .io_csrCtrl_eentry                               (cpuClockingArea_csr_io_ctrl_eentry[31:0]                                    ), //i
    .io_csrCtrl_tlbrentry                            (cpuClockingArea_csr_io_ctrl_tlbrentry[31:0]                                 ), //i
    .io_flush                                        (cpuClockingArea_rob_io_flush                                                ), //o
    .io_interrupt                                    (cpuClockingArea_csr_io_interrupt                                            ), //i
    .io_redirectPC                                   (cpuClockingArea_rob_io_redirectPC[31:0]                                     ), //o
    .io_commitROBEntries_0_pc                        (cpuClockingArea_rob_io_commitROBEntries_0_pc[31:0]                          ), //o
    .io_commitROBEntries_0_ard                       (cpuClockingArea_rob_io_commitROBEntries_0_ard[4:0]                          ), //o
    .io_commitROBEntries_0_prd                       (cpuClockingArea_rob_io_commitROBEntries_0_prd[5:0]                          ), //o
    .io_commitROBEntries_0_pprd                      (cpuClockingArea_rob_io_commitROBEntries_0_pprd[5:0]                         ), //o
    .io_commitROBEntries_0_specialOp                 (cpuClockingArea_rob_io_commitROBEntries_0_specialOp[3:0]                    ), //o
    .io_commitROBEntries_0_isComplete                (cpuClockingArea_rob_io_commitROBEntries_0_isComplete                        ), //o
    .io_commitROBEntries_0_branchResult_targetPC     (cpuClockingArea_rob_io_commitROBEntries_0_branchResult_targetPC[31:0]       ), //o
    .io_commitROBEntries_0_branchResult_branchResult (cpuClockingArea_rob_io_commitROBEntries_0_branchResult_branchResult         ), //o
    .io_commitROBEntries_0_branchResult_predictFail  (cpuClockingArea_rob_io_commitROBEntries_0_branchResult_predictFail          ), //o
    .io_commitROBEntries_0_exceptionInfo_exception   (cpuClockingArea_rob_io_commitROBEntries_0_exceptionInfo_exception           ), //o
    .io_commitROBEntries_0_exceptionInfo_eCode       (cpuClockingArea_rob_io_commitROBEntries_0_exceptionInfo_eCode[5:0]          ), //o
    .io_commitROBEntries_0_exceptionInfo_eSubCode    (cpuClockingArea_rob_io_commitROBEntries_0_exceptionInfo_eSubCode            ), //o
    .io_commitROBEntries_0_valid                     (cpuClockingArea_rob_io_commitROBEntries_0_valid                             ), //o
    .io_commitROBEntries_1_pc                        (cpuClockingArea_rob_io_commitROBEntries_1_pc[31:0]                          ), //o
    .io_commitROBEntries_1_ard                       (cpuClockingArea_rob_io_commitROBEntries_1_ard[4:0]                          ), //o
    .io_commitROBEntries_1_prd                       (cpuClockingArea_rob_io_commitROBEntries_1_prd[5:0]                          ), //o
    .io_commitROBEntries_1_pprd                      (cpuClockingArea_rob_io_commitROBEntries_1_pprd[5:0]                         ), //o
    .io_commitROBEntries_1_specialOp                 (cpuClockingArea_rob_io_commitROBEntries_1_specialOp[3:0]                    ), //o
    .io_commitROBEntries_1_isComplete                (cpuClockingArea_rob_io_commitROBEntries_1_isComplete                        ), //o
    .io_commitROBEntries_1_branchResult_targetPC     (cpuClockingArea_rob_io_commitROBEntries_1_branchResult_targetPC[31:0]       ), //o
    .io_commitROBEntries_1_branchResult_branchResult (cpuClockingArea_rob_io_commitROBEntries_1_branchResult_branchResult         ), //o
    .io_commitROBEntries_1_branchResult_predictFail  (cpuClockingArea_rob_io_commitROBEntries_1_branchResult_predictFail          ), //o
    .io_commitROBEntries_1_exceptionInfo_exception   (cpuClockingArea_rob_io_commitROBEntries_1_exceptionInfo_exception           ), //o
    .io_commitROBEntries_1_exceptionInfo_eCode       (cpuClockingArea_rob_io_commitROBEntries_1_exceptionInfo_eCode[5:0]          ), //o
    .io_commitROBEntries_1_exceptionInfo_eSubCode    (cpuClockingArea_rob_io_commitROBEntries_1_exceptionInfo_eSubCode            ), //o
    .io_commitROBEntries_1_valid                     (cpuClockingArea_rob_io_commitROBEntries_1_valid                             ), //o
    .io_commitROBEntries_2_pc                        (cpuClockingArea_rob_io_commitROBEntries_2_pc[31:0]                          ), //o
    .io_commitROBEntries_2_ard                       (cpuClockingArea_rob_io_commitROBEntries_2_ard[4:0]                          ), //o
    .io_commitROBEntries_2_prd                       (cpuClockingArea_rob_io_commitROBEntries_2_prd[5:0]                          ), //o
    .io_commitROBEntries_2_pprd                      (cpuClockingArea_rob_io_commitROBEntries_2_pprd[5:0]                         ), //o
    .io_commitROBEntries_2_specialOp                 (cpuClockingArea_rob_io_commitROBEntries_2_specialOp[3:0]                    ), //o
    .io_commitROBEntries_2_isComplete                (cpuClockingArea_rob_io_commitROBEntries_2_isComplete                        ), //o
    .io_commitROBEntries_2_branchResult_targetPC     (cpuClockingArea_rob_io_commitROBEntries_2_branchResult_targetPC[31:0]       ), //o
    .io_commitROBEntries_2_branchResult_branchResult (cpuClockingArea_rob_io_commitROBEntries_2_branchResult_branchResult         ), //o
    .io_commitROBEntries_2_branchResult_predictFail  (cpuClockingArea_rob_io_commitROBEntries_2_branchResult_predictFail          ), //o
    .io_commitROBEntries_2_exceptionInfo_exception   (cpuClockingArea_rob_io_commitROBEntries_2_exceptionInfo_exception           ), //o
    .io_commitROBEntries_2_exceptionInfo_eCode       (cpuClockingArea_rob_io_commitROBEntries_2_exceptionInfo_eCode[5:0]          ), //o
    .io_commitROBEntries_2_exceptionInfo_eSubCode    (cpuClockingArea_rob_io_commitROBEntries_2_exceptionInfo_eSubCode            ), //o
    .io_commitROBEntries_2_valid                     (cpuClockingArea_rob_io_commitROBEntries_2_valid                             ), //o
    .io_commitROBEntries_3_pc                        (cpuClockingArea_rob_io_commitROBEntries_3_pc[31:0]                          ), //o
    .io_commitROBEntries_3_ard                       (cpuClockingArea_rob_io_commitROBEntries_3_ard[4:0]                          ), //o
    .io_commitROBEntries_3_prd                       (cpuClockingArea_rob_io_commitROBEntries_3_prd[5:0]                          ), //o
    .io_commitROBEntries_3_pprd                      (cpuClockingArea_rob_io_commitROBEntries_3_pprd[5:0]                         ), //o
    .io_commitROBEntries_3_specialOp                 (cpuClockingArea_rob_io_commitROBEntries_3_specialOp[3:0]                    ), //o
    .io_commitROBEntries_3_isComplete                (cpuClockingArea_rob_io_commitROBEntries_3_isComplete                        ), //o
    .io_commitROBEntries_3_branchResult_targetPC     (cpuClockingArea_rob_io_commitROBEntries_3_branchResult_targetPC[31:0]       ), //o
    .io_commitROBEntries_3_branchResult_branchResult (cpuClockingArea_rob_io_commitROBEntries_3_branchResult_branchResult         ), //o
    .io_commitROBEntries_3_branchResult_predictFail  (cpuClockingArea_rob_io_commitROBEntries_3_branchResult_predictFail          ), //o
    .io_commitROBEntries_3_exceptionInfo_exception   (cpuClockingArea_rob_io_commitROBEntries_3_exceptionInfo_exception           ), //o
    .io_commitROBEntries_3_exceptionInfo_eCode       (cpuClockingArea_rob_io_commitROBEntries_3_exceptionInfo_eCode[5:0]          ), //o
    .io_commitROBEntries_3_exceptionInfo_eSubCode    (cpuClockingArea_rob_io_commitROBEntries_3_exceptionInfo_eSubCode            ), //o
    .io_commitROBEntries_3_valid                     (cpuClockingArea_rob_io_commitROBEntries_3_valid                             ), //o
    .io_commitROBEntries_4_pc                        (cpuClockingArea_rob_io_commitROBEntries_4_pc[31:0]                          ), //o
    .io_commitROBEntries_4_ard                       (cpuClockingArea_rob_io_commitROBEntries_4_ard[4:0]                          ), //o
    .io_commitROBEntries_4_prd                       (cpuClockingArea_rob_io_commitROBEntries_4_prd[5:0]                          ), //o
    .io_commitROBEntries_4_pprd                      (cpuClockingArea_rob_io_commitROBEntries_4_pprd[5:0]                         ), //o
    .io_commitROBEntries_4_specialOp                 (cpuClockingArea_rob_io_commitROBEntries_4_specialOp[3:0]                    ), //o
    .io_commitROBEntries_4_isComplete                (cpuClockingArea_rob_io_commitROBEntries_4_isComplete                        ), //o
    .io_commitROBEntries_4_branchResult_targetPC     (cpuClockingArea_rob_io_commitROBEntries_4_branchResult_targetPC[31:0]       ), //o
    .io_commitROBEntries_4_branchResult_branchResult (cpuClockingArea_rob_io_commitROBEntries_4_branchResult_branchResult         ), //o
    .io_commitROBEntries_4_branchResult_predictFail  (cpuClockingArea_rob_io_commitROBEntries_4_branchResult_predictFail          ), //o
    .io_commitROBEntries_4_exceptionInfo_exception   (cpuClockingArea_rob_io_commitROBEntries_4_exceptionInfo_exception           ), //o
    .io_commitROBEntries_4_exceptionInfo_eCode       (cpuClockingArea_rob_io_commitROBEntries_4_exceptionInfo_eCode[5:0]          ), //o
    .io_commitROBEntries_4_exceptionInfo_eSubCode    (cpuClockingArea_rob_io_commitROBEntries_4_exceptionInfo_eSubCode            ), //o
    .io_commitROBEntries_4_valid                     (cpuClockingArea_rob_io_commitROBEntries_4_valid                             ), //o
    .aclk                                            (aclk                                                                        ), //i
    .aresetn                                         (aresetn                                                                     )  //i
  );
  CSR cpuClockingArea_csr (
    .io_extInt                       (intrpt[7:0]                                                    ), //i
    .io_interrupt                    (cpuClockingArea_csr_io_interrupt                               ), //o
    ._zz_when_Cache_l83              (cpuClockingArea_csr__zz_when_Cache_l83[1:0]                    ), //o
    .io_counter_id                   (cpuClockingArea_csr_io_counter_id[31:0]                        ), //o
    .io_counter_value                (cpuClockingArea_csr_io_counter_value[63:0]                     ), //o
    .io_swRead_value                 (cpuClockingArea_csr_io_swRead_value[31:0]                      ), //o
    .io_swRead_address               (cpuClockingArea_areaFlushReset_roALU0_io_csr_address[13:0]     ), //i
    .io_swWrite_value                (cpuClockingArea_areaFlushReset_fuALU0_io_csrWrite_value[31:0]  ), //i
    .io_swWrite_address              (cpuClockingArea_areaFlushReset_fuALU0_io_csrWrite_address[13:0]), //i
    .io_swWrite_wen                  (cpuClockingArea_areaFlushReset_fuALU0_io_csrWrite_wen          ), //i
    .io_llBitComm_actualAddr         (cpuClockingArea_csr_io_llBitComm_actualAddr[31:0]              ), //o
    .io_llBitComm_toUpdateAddr       (cpuClockingArea_fuLSU_io_llBitComm_toUpdateAddr[31:0]          ), //i
    .io_llBitComm_wen                (cpuClockingArea_fuLSU_io_llBitComm_wen                         ), //i
    ._zz_scMatchHit                  (cpuClockingArea_csr__zz_scMatchHit                             ), //o
    .io_badvICache_vaddr             (cpuClockingArea_iCache_io_badv_vaddr[31:0]                     ), //i
    .io_badvICache_wen               (cpuClockingArea_iCache_io_badv_wen                             ), //i
    .io_badvDCache_robIdx            (cpuClockingArea_fuLSU_io_badv_robIdx[4:0]                      ), //i
    .io_badvDCache_vaddr             (cpuClockingArea_fuLSU_io_badv_vaddr[31:0]                      ), //i
    .io_badvDCache_wen               (cpuClockingArea_fuLSU_io_badv_wen                              ), //i
    .io_tlbCSRInfo_asid              (cpuClockingArea_csr_io_tlbCSRInfo_asid[9:0]                    ), //o
    ._zz_io_iCacheReq_pageInfo_plv   (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_plv[1:0]         ), //o
    ._zz_when_TLB_l177               (cpuClockingArea_csr__zz_when_TLB_l177                          ), //o
    ._zz_when_TLB_l177_1             (cpuClockingArea_csr__zz_when_TLB_l177_1                        ), //o
    ._zz_io_iCacheReq_pageInfo_mat   (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_mat[1:0]         ), //o
    ._zz_io_dCacheReq_pageInfo_mat   (cpuClockingArea_csr__zz_io_dCacheReq_pageInfo_mat[1:0]         ), //o
    ._zz_when_TLB_l178               (cpuClockingArea_csr__zz_when_TLB_l178                          ), //o
    ._zz_when_TLB_l178_1             (cpuClockingArea_csr__zz_when_TLB_l178_1                        ), //o
    ._zz_io_iCacheReq_pageInfo_mat_1 (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_mat_1[1:0]       ), //o
    ._zz_io_iCacheReq_pageInfo_ppn   (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_ppn[2:0]         ), //o
    ._zz_when_TLB_l178_2             (cpuClockingArea_csr__zz_when_TLB_l178_2[2:0]                   ), //o
    ._zz_when_TLB_l185               (cpuClockingArea_csr__zz_when_TLB_l185                          ), //o
    ._zz_when_TLB_l185_1             (cpuClockingArea_csr__zz_when_TLB_l185_1                        ), //o
    ._zz_io_iCacheReq_pageInfo_mat_2 (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_mat_2[1:0]       ), //o
    ._zz_io_iCacheReq_pageInfo_ppn_1 (cpuClockingArea_csr__zz_io_iCacheReq_pageInfo_ppn_1[2:0]       ), //o
    ._zz_when_TLB_l185_2             (cpuClockingArea_csr__zz_when_TLB_l185_2[2:0]                   ), //o
    ._zz_entryToFill_e               (cpuClockingArea_csr__zz_entryToFill_e[5:0]                     ), //o
    ._zz_io_csrWrite_asid            (cpuClockingArea_csr__zz_io_csrWrite_asid[1:0]                  ), //o
    ._zz_io_swRead_value             (cpuClockingArea_csr__zz_io_swRead_value[21:0]                  ), //o
    ._zz_entryToFill_ps              (cpuClockingArea_csr__zz_entryToFill_ps[5:0]                    ), //o
    ._zz_io_swRead_value_1           (cpuClockingArea_csr__zz_io_swRead_value_1                      ), //o
    ._zz_entryToFill_e_1             (cpuClockingArea_csr__zz_entryToFill_e_1                        ), //o
    ._zz_entryToFill_vppn            (cpuClockingArea_csr__zz_entryToFill_vppn[18:0]                 ), //o
    ._zz_entryToFill_pp0_v           (cpuClockingArea_csr__zz_entryToFill_pp0_v                      ), //o
    ._zz_entryToFill_pp0_d           (cpuClockingArea_csr__zz_entryToFill_pp0_d                      ), //o
    ._zz_entryToFill_pp0_plv         (cpuClockingArea_csr__zz_entryToFill_pp0_plv[1:0]               ), //o
    ._zz_entryToFill_pp0_mat         (cpuClockingArea_csr__zz_entryToFill_pp0_mat[1:0]               ), //o
    ._zz_entryToFill_g               (cpuClockingArea_csr__zz_entryToFill_g                          ), //o
    ._zz_entryToFill_pp0_ppn         (cpuClockingArea_csr__zz_entryToFill_pp0_ppn[19:0]              ), //o
    ._zz_entryToFill_pp1_v           (cpuClockingArea_csr__zz_entryToFill_pp1_v                      ), //o
    ._zz_entryToFill_pp1_d           (cpuClockingArea_csr__zz_entryToFill_pp1_d                      ), //o
    ._zz_entryToFill_pp1_plv         (cpuClockingArea_csr__zz_entryToFill_pp1_plv[1:0]               ), //o
    ._zz_entryToFill_pp1_mat         (cpuClockingArea_csr__zz_entryToFill_pp1_mat[1:0]               ), //o
    ._zz_entryToFill_g_1             (cpuClockingArea_csr__zz_entryToFill_g_1                        ), //o
    ._zz_entryToFill_pp1_ppn         (cpuClockingArea_csr__zz_entryToFill_pp1_ppn[19:0]              ), //o
    ._zz_io_swRead_value_2           (cpuClockingArea_tlb__zz_io_swRead_value_2[1:0]                 ), //i
    ._zz_io_swRead_value_3           (cpuClockingArea_tlb__zz_io_swRead_value_3[21:0]                ), //i
    ._zz_io_swRead_value_4           (cpuClockingArea_tlb__zz_io_swRead_value_4[5:0]                 ), //i
    ._zz_io_swRead_value_5           (cpuClockingArea_tlb__zz_io_swRead_value_5                      ), //i
    ._zz_io_swRead_value_6           (cpuClockingArea_tlb__zz_io_swRead_value_6                      ), //i
    ._zz_io_swRead_value_7           (cpuClockingArea_tlb__zz_io_swRead_value_7[12:0]                ), //i
    ._zz_io_swRead_value_8           (cpuClockingArea_tlb__zz_io_swRead_value_8[18:0]                ), //i
    ._zz_io_swRead_value_9           (cpuClockingArea_tlb__zz_io_swRead_value_9                      ), //i
    ._zz_io_swRead_value_10          (cpuClockingArea_tlb__zz_io_swRead_value_10                     ), //i
    ._zz_io_swRead_value_11          (cpuClockingArea_tlb__zz_io_swRead_value_11[1:0]                ), //i
    ._zz_io_swRead_value_12          (cpuClockingArea_tlb__zz_io_swRead_value_12[1:0]                ), //i
    ._zz_io_swRead_value_13          (cpuClockingArea_tlb__zz_io_swRead_value_13                     ), //i
    ._zz_io_swRead_value_14          (cpuClockingArea_tlb__zz_io_swRead_value_14                     ), //i
    ._zz_io_swRead_value_15          (cpuClockingArea_tlb__zz_io_swRead_value_15[19:0]               ), //i
    ._zz_io_swRead_value_16          (cpuClockingArea_tlb__zz_io_swRead_value_16[3:0]                ), //i
    ._zz_io_swRead_value_17          (cpuClockingArea_tlb__zz_io_swRead_value_17                     ), //i
    ._zz_io_swRead_value_18          (cpuClockingArea_tlb__zz_io_swRead_value_18                     ), //i
    ._zz_io_swRead_value_19          (cpuClockingArea_tlb__zz_io_swRead_value_19[1:0]                ), //i
    ._zz_io_swRead_value_20          (cpuClockingArea_tlb__zz_io_swRead_value_20[1:0]                ), //i
    ._zz_io_swRead_value_21          (cpuClockingArea_tlb__zz_io_swRead_value_21                     ), //i
    ._zz_io_swRead_value_22          (cpuClockingArea_tlb__zz_io_swRead_value_22                     ), //i
    ._zz_io_swRead_value_23          (cpuClockingArea_tlb__zz_io_swRead_value_23[19:0]               ), //i
    ._zz_io_swRead_value_24          (cpuClockingArea_tlb__zz_io_swRead_value_24[3:0]                ), //i
    .io_tlbCSRWrite_asid             (cpuClockingArea_tlb_io_csrWrite_asid[9:0]                      ), //i
    .io_tlbCSRWrite_idxWen           (cpuClockingArea_tlb_io_csrWrite_idxWen                         ), //i
    .io_tlbCSRWrite_entryWen         (cpuClockingArea_tlb_io_csrWrite_entryWen                       ), //i
    .io_ctrl_llBitUpdate             (cpuClockingArea_rob_io_csrCtrl_llBitUpdate                     ), //i
    .io_ctrl_writeCSR                (cpuClockingArea_rob_io_csrCtrl_writeCSR                        ), //i
    .io_ctrl_ertn                    (cpuClockingArea_rob_io_csrCtrl_ertn                            ), //i
    .io_ctrl_normalException         (cpuClockingArea_rob_io_csrCtrl_normalException                 ), //i
    .io_ctrl_tlbrException           (cpuClockingArea_rob_io_csrCtrl_tlbrException                   ), //i
    .io_ctrl_epc                     (cpuClockingArea_rob_io_csrCtrl_epc[31:0]                       ), //i
    .io_ctrl_eROBIdx                 (cpuClockingArea_rob_io_csrCtrl_eROBIdx[4:0]                    ), //i
    .io_ctrl_eCode                   (cpuClockingArea_rob_io_csrCtrl_eCode[5:0]                      ), //i
    .io_ctrl_eSubCode                (cpuClockingArea_rob_io_csrCtrl_eSubCode                        ), //i
    .io_ctrl_era                     (cpuClockingArea_csr_io_ctrl_era[31:0]                          ), //o
    .io_ctrl_eentry                  (cpuClockingArea_csr_io_ctrl_eentry[31:0]                       ), //o
    .io_ctrl_tlbrentry               (cpuClockingArea_csr_io_ctrl_tlbrentry[31:0]                    ), //o
    .io_flush                        (cpuClockingArea_rob_io_flush                                   ), //i
    .io_diffCSRBundle_crmd           (cpuClockingArea_csr_io_diffCSRBundle_crmd[31:0]                ), //o
    .io_diffCSRBundle_prmd           (cpuClockingArea_csr_io_diffCSRBundle_prmd[31:0]                ), //o
    .io_diffCSRBundle_ecfg           (cpuClockingArea_csr_io_diffCSRBundle_ecfg[31:0]                ), //o
    .io_diffCSRBundle_estat          (cpuClockingArea_csr_io_diffCSRBundle_estat[31:0]               ), //o
    .io_diffCSRBundle_era            (cpuClockingArea_csr_io_diffCSRBundle_era[31:0]                 ), //o
    .io_diffCSRBundle_badv           (cpuClockingArea_csr_io_diffCSRBundle_badv[31:0]                ), //o
    .io_diffCSRBundle_eentry         (cpuClockingArea_csr_io_diffCSRBundle_eentry[31:0]              ), //o
    .io_diffCSRBundle_tlbidx         (cpuClockingArea_csr_io_diffCSRBundle_tlbidx[31:0]              ), //o
    .io_diffCSRBundle_tlbehi         (cpuClockingArea_csr_io_diffCSRBundle_tlbehi[31:0]              ), //o
    .io_diffCSRBundle_tlbelo0        (cpuClockingArea_csr_io_diffCSRBundle_tlbelo0[31:0]             ), //o
    .io_diffCSRBundle_tlbelo1        (cpuClockingArea_csr_io_diffCSRBundle_tlbelo1[31:0]             ), //o
    .io_diffCSRBundle_asid           (cpuClockingArea_csr_io_diffCSRBundle_asid[31:0]                ), //o
    .io_diffCSRBundle_pgdl           (cpuClockingArea_csr_io_diffCSRBundle_pgdl[31:0]                ), //o
    .io_diffCSRBundle_pgdh           (cpuClockingArea_csr_io_diffCSRBundle_pgdh[31:0]                ), //o
    .io_diffCSRBundle_save0          (cpuClockingArea_csr_io_diffCSRBundle_save0[31:0]               ), //o
    .io_diffCSRBundle_save1          (cpuClockingArea_csr_io_diffCSRBundle_save1[31:0]               ), //o
    .io_diffCSRBundle_save2          (cpuClockingArea_csr_io_diffCSRBundle_save2[31:0]               ), //o
    .io_diffCSRBundle_save3          (cpuClockingArea_csr_io_diffCSRBundle_save3[31:0]               ), //o
    .io_diffCSRBundle_tid            (cpuClockingArea_csr_io_diffCSRBundle_tid[31:0]                 ), //o
    .io_diffCSRBundle_tcfg           (cpuClockingArea_csr_io_diffCSRBundle_tcfg[31:0]                ), //o
    .io_diffCSRBundle_tval           (cpuClockingArea_csr_io_diffCSRBundle_tval[31:0]                ), //o
    .io_diffCSRBundle_ticlr          (cpuClockingArea_csr_io_diffCSRBundle_ticlr[31:0]               ), //o
    .io_diffCSRBundle_llbctl         (cpuClockingArea_csr_io_diffCSRBundle_llbctl[31:0]              ), //o
    .io_diffCSRBundle_tlbrentry      (cpuClockingArea_csr_io_diffCSRBundle_tlbrentry[31:0]           ), //o
    .io_diffCSRBundle_dmw0           (cpuClockingArea_csr_io_diffCSRBundle_dmw0[31:0]                ), //o
    .io_diffCSRBundle_dmw1           (cpuClockingArea_csr_io_diffCSRBundle_dmw1[31:0]                ), //o
    .aclk                            (aclk                                                           ), //i
    .aresetn                         (aresetn                                                        )  //i
  );
  InstrQueue cpuClockingArea_areaFlushReset_instQueue (
    .io_in_allowMask                         (cpuClockingArea_areaFlushReset_instQueue_io_in_allowMask[1:0]                    ), //o
    .io_in_availMask                         (cpuClockingArea_iCache_io_output_availMask[1:0]                                  ), //i
    .io_in_info_0_inst                       (cpuClockingArea_iCache_io_output_info_0_inst[31:0]                               ), //i
    .io_in_info_0_branchInfo_predictPC       (cpuClockingArea_iCache_io_output_info_0_branchInfo_predictPC[31:0]               ), //i
    .io_in_info_0_branchInfo_predictResult   (cpuClockingArea_iCache_io_output_info_0_branchInfo_predictResult                 ), //i
    .io_in_info_0_exceptionInfo_exception    (cpuClockingArea_iCache_io_output_info_0_exceptionInfo_exception                  ), //i
    .io_in_info_0_exceptionInfo_eCode        (cpuClockingArea_iCache_io_output_info_0_exceptionInfo_eCode[5:0]                 ), //i
    .io_in_info_0_exceptionInfo_eSubCode     (cpuClockingArea_iCache_io_output_info_0_exceptionInfo_eSubCode                   ), //i
    .io_in_info_0_pc                         (cpuClockingArea_iCache_io_output_info_0_pc[31:0]                                 ), //i
    .io_in_info_1_inst                       (cpuClockingArea_iCache_io_output_info_1_inst[31:0]                               ), //i
    .io_in_info_1_branchInfo_predictPC       (cpuClockingArea_iCache_io_output_info_1_branchInfo_predictPC[31:0]               ), //i
    .io_in_info_1_branchInfo_predictResult   (cpuClockingArea_iCache_io_output_info_1_branchInfo_predictResult                 ), //i
    .io_in_info_1_exceptionInfo_exception    (cpuClockingArea_iCache_io_output_info_1_exceptionInfo_exception                  ), //i
    .io_in_info_1_exceptionInfo_eCode        (cpuClockingArea_iCache_io_output_info_1_exceptionInfo_eCode[5:0]                 ), //i
    .io_in_info_1_exceptionInfo_eSubCode     (cpuClockingArea_iCache_io_output_info_1_exceptionInfo_eSubCode                   ), //i
    .io_in_info_1_pc                         (cpuClockingArea_iCache_io_output_info_1_pc[31:0]                                 ), //i
    .io_out_allowMask                        (cpuClockingArea_areaFlushReset_dispatcher_io_input_allowMask[1:0]                ), //i
    .io_out_availMask                        (cpuClockingArea_areaFlushReset_instQueue_io_out_availMask[1:0]                   ), //o
    .io_out_info_0_inst                      (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_inst[31:0]                ), //o
    .io_out_info_0_branchInfo_predictPC      (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_branchInfo_predictPC[31:0]), //o
    .io_out_info_0_branchInfo_predictResult  (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_branchInfo_predictResult  ), //o
    .io_out_info_0_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_exceptionInfo_exception   ), //o
    .io_out_info_0_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_exceptionInfo_eCode[5:0]  ), //o
    .io_out_info_0_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_exceptionInfo_eSubCode    ), //o
    .io_out_info_0_pc                        (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_pc[31:0]                  ), //o
    .io_out_info_1_inst                      (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_inst[31:0]                ), //o
    .io_out_info_1_branchInfo_predictPC      (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_branchInfo_predictPC[31:0]), //o
    .io_out_info_1_branchInfo_predictResult  (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_branchInfo_predictResult  ), //o
    .io_out_info_1_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_exceptionInfo_exception   ), //o
    .io_out_info_1_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_exceptionInfo_eCode[5:0]  ), //o
    .io_out_info_1_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_exceptionInfo_eSubCode    ), //o
    .io_out_info_1_pc                        (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_pc[31:0]                  ), //o
    .io_out_dispatchInfo_0_fuType            (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_fuType[2:0]       ), //o
    .io_out_dispatchInfo_0_ard               (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_ard[4:0]          ), //o
    .io_out_dispatchInfo_0_asrc_0            (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_asrc_0[4:0]       ), //o
    .io_out_dispatchInfo_0_asrc_1            (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_asrc_1[4:0]       ), //o
    .io_out_dispatchInfo_1_fuType            (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_fuType[2:0]       ), //o
    .io_out_dispatchInfo_1_ard               (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_ard[4:0]          ), //o
    .io_out_dispatchInfo_1_asrc_0            (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_asrc_0[4:0]       ), //o
    .io_out_dispatchInfo_1_asrc_1            (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_asrc_1[4:0]       ), //o
    .aclk                                    (aclk                                                                             ), //i
    .cpuClockingArea_areaFlushReset_newReset (cpuClockingArea_areaFlushReset_newReset                                          )  //i
  );
  Dispatcher cpuClockingArea_areaFlushReset_dispatcher (
    .io_input_allowMask                          (cpuClockingArea_areaFlushReset_dispatcher_io_input_allowMask[1:0]                      ), //o
    .io_input_availMask                          (cpuClockingArea_areaFlushReset_instQueue_io_out_availMask[1:0]                         ), //i
    .io_input_info_0_inst                        (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_inst[31:0]                      ), //i
    .io_input_info_0_branchInfo_predictPC        (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_branchInfo_predictPC[31:0]      ), //i
    .io_input_info_0_branchInfo_predictResult    (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_branchInfo_predictResult        ), //i
    .io_input_info_0_exceptionInfo_exception     (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_exceptionInfo_exception         ), //i
    .io_input_info_0_exceptionInfo_eCode         (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_exceptionInfo_eCode[5:0]        ), //i
    .io_input_info_0_exceptionInfo_eSubCode      (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_exceptionInfo_eSubCode          ), //i
    .io_input_info_0_pc                          (cpuClockingArea_areaFlushReset_instQueue_io_out_info_0_pc[31:0]                        ), //i
    .io_input_info_1_inst                        (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_inst[31:0]                      ), //i
    .io_input_info_1_branchInfo_predictPC        (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_branchInfo_predictPC[31:0]      ), //i
    .io_input_info_1_branchInfo_predictResult    (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_branchInfo_predictResult        ), //i
    .io_input_info_1_exceptionInfo_exception     (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_exceptionInfo_exception         ), //i
    .io_input_info_1_exceptionInfo_eCode         (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_exceptionInfo_eCode[5:0]        ), //i
    .io_input_info_1_exceptionInfo_eSubCode      (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_exceptionInfo_eSubCode          ), //i
    .io_input_info_1_pc                          (cpuClockingArea_areaFlushReset_instQueue_io_out_info_1_pc[31:0]                        ), //i
    .io_input_dispatchInfo_0_fuType              (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_fuType[2:0]             ), //i
    .io_input_dispatchInfo_0_ard                 (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_ard[4:0]                ), //i
    .io_input_dispatchInfo_0_asrc_0              (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_asrc_0[4:0]             ), //i
    .io_input_dispatchInfo_0_asrc_1              (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_0_asrc_1[4:0]             ), //i
    .io_input_dispatchInfo_1_fuType              (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_fuType[2:0]             ), //i
    .io_input_dispatchInfo_1_ard                 (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_ard[4:0]                ), //i
    .io_input_dispatchInfo_1_asrc_0              (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_asrc_0[4:0]             ), //i
    .io_input_dispatchInfo_1_asrc_1              (cpuClockingArea_areaFlushReset_instQueue_io_out_dispatchInfo_1_asrc_1[4:0]             ), //i
    .io_aluHasCSRInst_0                          (cpuClockingArea_areaFlushReset_issueQueueALU0_io_csrInQueue                            ), //i
    .io_aluHasCSRInst_1                          (cpuClockingArea_areaFlushReset_issueQueueALU1_io_csrInQueue                            ), //i
    .io_rob_allowMask                            (cpuClockingArea_areaFlushReset_dispatcher_io_rob_allowMask[1:0]                        ), //o
    .io_rob_availMask                            (cpuClockingArea_rob_io_dispatch_availMask[1:0]                                         ), //i
    .io_rob_robIdx_0                             (cpuClockingArea_rob_io_dispatch_robIdx_0[4:0]                                          ), //i
    .io_rob_robIdx_1                             (cpuClockingArea_rob_io_dispatch_robIdx_1[4:0]                                          ), //i
    .io_rob_pc_0                                 (cpuClockingArea_areaFlushReset_dispatcher_io_rob_pc_0[31:0]                            ), //o
    .io_rob_pc_1                                 (cpuClockingArea_areaFlushReset_dispatcher_io_rob_pc_1[31:0]                            ), //o
    .io_rob_ard_0                                (cpuClockingArea_areaFlushReset_dispatcher_io_rob_ard_0[4:0]                            ), //o
    .io_rob_ard_1                                (cpuClockingArea_areaFlushReset_dispatcher_io_rob_ard_1[4:0]                            ), //o
    .io_rob_prd_0                                (cpuClockingArea_areaFlushReset_dispatcher_io_rob_prd_0[5:0]                            ), //o
    .io_rob_prd_1                                (cpuClockingArea_areaFlushReset_dispatcher_io_rob_prd_1[5:0]                            ), //o
    .io_rob_pprd_0                               (cpuClockingArea_areaFlushReset_dispatcher_io_rob_pprd_0[5:0]                           ), //o
    .io_rob_pprd_1                               (cpuClockingArea_areaFlushReset_dispatcher_io_rob_pprd_1[5:0]                           ), //o
    .io_rob_specialOp_0                          (cpuClockingArea_areaFlushReset_dispatcher_io_rob_specialOp_0[3:0]                      ), //o
    .io_rob_specialOp_1                          (cpuClockingArea_areaFlushReset_dispatcher_io_rob_specialOp_1[3:0]                      ), //o
    .io_sratWrite_0_ard                          (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_0_ard[4:0]                      ), //o
    .io_sratWrite_0_prd                          (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_0_prd[5:0]                      ), //o
    .io_sratWrite_0_wen                          (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_0_wen                           ), //o
    .io_sratWrite_1_ard                          (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_1_ard[4:0]                      ), //o
    .io_sratWrite_1_prd                          (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_1_prd[5:0]                      ), //o
    .io_sratWrite_1_wen                          (cpuClockingArea_areaFlushReset_dispatcher_io_sratWrite_1_wen                           ), //o
    .io_sratReadSrc_0_0_ard                      (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_0_0_ard[4:0]                  ), //o
    .io_sratReadSrc_0_0_prd                      (cpuClockingArea_sRAT_io_srcReadPort_0_0_prd[5:0]                                       ), //i
    .io_sratReadSrc_0_0_valid                    (cpuClockingArea_sRAT_io_srcReadPort_0_0_valid                                          ), //i
    .io_sratReadSrc_0_1_ard                      (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_0_1_ard[4:0]                  ), //o
    .io_sratReadSrc_0_1_prd                      (cpuClockingArea_sRAT_io_srcReadPort_0_1_prd[5:0]                                       ), //i
    .io_sratReadSrc_0_1_valid                    (cpuClockingArea_sRAT_io_srcReadPort_0_1_valid                                          ), //i
    .io_sratReadSrc_1_0_ard                      (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_1_0_ard[4:0]                  ), //o
    .io_sratReadSrc_1_0_prd                      (cpuClockingArea_sRAT_io_srcReadPort_1_0_prd[5:0]                                       ), //i
    .io_sratReadSrc_1_0_valid                    (cpuClockingArea_sRAT_io_srcReadPort_1_0_valid                                          ), //i
    .io_sratReadSrc_1_1_ard                      (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadSrc_1_1_ard[4:0]                  ), //o
    .io_sratReadSrc_1_1_prd                      (cpuClockingArea_sRAT_io_srcReadPort_1_1_prd[5:0]                                       ), //i
    .io_sratReadSrc_1_1_valid                    (cpuClockingArea_sRAT_io_srcReadPort_1_1_valid                                          ), //i
    .io_sratReadPPRD_0_ard                       (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadPPRD_0_ard[4:0]                   ), //o
    .io_sratReadPPRD_0_prd                       (cpuClockingArea_sRAT_io_prevPRDReadPort_0_prd[5:0]                                     ), //i
    .io_sratReadPPRD_0_valid                     (cpuClockingArea_sRAT_io_prevPRDReadPort_0_valid                                        ), //i
    .io_sratReadPPRD_1_ard                       (cpuClockingArea_areaFlushReset_dispatcher_io_sratReadPPRD_1_ard[4:0]                   ), //o
    .io_sratReadPPRD_1_prd                       (cpuClockingArea_sRAT_io_prevPRDReadPort_1_prd[5:0]                                     ), //i
    .io_sratReadPPRD_1_valid                     (cpuClockingArea_sRAT_io_prevPRDReadPort_1_valid                                        ), //i
    .io_freelist_disPatchNum                     (cpuClockingArea_areaFlushReset_dispatcher_io_freelist_disPatchNum[1:0]                 ), //o
    .io_freelist_availMask                       (cpuClockingArea_freeList_io_dispatch_availMask[1:0]                                    ), //i
    .io_freelist_prfIdx_0                        (cpuClockingArea_freeList_io_dispatch_prfIdx_0[5:0]                                     ), //i
    .io_freelist_prfIdx_1                        (cpuClockingArea_freeList_io_dispatch_prfIdx_1[5:0]                                     ), //i
    ._zz_when_Decoder_l40                        (cpuClockingArea_csr__zz_when_Cache_l83[1:0]                                            ), //i
    .io_alu0IQ_valid                             (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_valid                              ), //o
    .io_alu0IQ_ready                             (cpuClockingArea_areaFlushReset_issueQueueALU0_io_input_ready                           ), //i
    .io_alu0IQ_payload_robIdx                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_robIdx[4:0]                ), //o
    .io_alu0IQ_payload_branchInfo_predictPC      (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_branchInfo_predictPC[31:0] ), //o
    .io_alu0IQ_payload_branchInfo_predictResult  (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_branchInfo_predictResult   ), //o
    .io_alu0IQ_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_exceptionInfo_exception    ), //o
    .io_alu0IQ_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_exceptionInfo_eCode[5:0]   ), //o
    .io_alu0IQ_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_exceptionInfo_eSubCode     ), //o
    .io_alu0IQ_payload_pc                        (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_pc[31:0]                   ), //o
    .io_alu0IQ_payload_prd                       (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_prd[5:0]                   ), //o
    .io_alu0IQ_payload_psrc_0                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_psrc_0[5:0]                ), //o
    .io_alu0IQ_payload_psrc_1                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_psrc_1[5:0]                ), //o
    .io_alu0IQ_payload_imm                       (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_imm[31:0]                  ), //o
    .io_alu0IQ_payload_uop_aluOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_uop_aluOp[3:0]             ), //o
    .io_alu0IQ_payload_uop_bruOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_uop_bruOp[1:0]             ), //o
    .io_alu0IQ_payload_uop_cruOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_uop_cruOp[1:0]             ), //o
    .io_alu0IQ_payload_roop_aluROOp              (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_roop_aluROOp[2:0]          ), //o
    .io_alu0IQ_payload_srcReady_0                (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_srcReady_0                 ), //o
    .io_alu0IQ_payload_srcReady_1                (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_srcReady_1                 ), //o
    .io_alu1IQ_valid                             (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_valid                              ), //o
    .io_alu1IQ_ready                             (cpuClockingArea_areaFlushReset_issueQueueALU1_io_input_ready                           ), //i
    .io_alu1IQ_payload_robIdx                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_robIdx[4:0]                ), //o
    .io_alu1IQ_payload_branchInfo_predictPC      (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_branchInfo_predictPC[31:0] ), //o
    .io_alu1IQ_payload_branchInfo_predictResult  (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_branchInfo_predictResult   ), //o
    .io_alu1IQ_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_exceptionInfo_exception    ), //o
    .io_alu1IQ_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_exceptionInfo_eCode[5:0]   ), //o
    .io_alu1IQ_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_exceptionInfo_eSubCode     ), //o
    .io_alu1IQ_payload_pc                        (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_pc[31:0]                   ), //o
    .io_alu1IQ_payload_prd                       (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_prd[5:0]                   ), //o
    .io_alu1IQ_payload_psrc_0                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_psrc_0[5:0]                ), //o
    .io_alu1IQ_payload_psrc_1                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_psrc_1[5:0]                ), //o
    .io_alu1IQ_payload_imm                       (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_imm[31:0]                  ), //o
    .io_alu1IQ_payload_uop_aluOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_uop_aluOp[3:0]             ), //o
    .io_alu1IQ_payload_uop_bruOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_uop_bruOp[1:0]             ), //o
    .io_alu1IQ_payload_roop_aluROOp              (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_roop_aluROOp[2:0]          ), //o
    .io_alu1IQ_payload_roop_cruROOp              (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_roop_cruROOp[1:0]          ), //o
    .io_alu1IQ_payload_srcReady_0                (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_srcReady_0                 ), //o
    .io_alu1IQ_payload_srcReady_1                (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_srcReady_1                 ), //o
    .io_muluIQ_valid                             (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_valid                              ), //o
    .io_muluIQ_ready                             (cpuClockingArea_areaFlushReset_issueQueueMULU_io_input_ready                           ), //i
    .io_muluIQ_payload_robIdx                    (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_robIdx[4:0]                ), //o
    .io_muluIQ_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_branchResult_targetPC[31:0]), //o
    .io_muluIQ_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_branchResult_branchResult  ), //o
    .io_muluIQ_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_branchResult_predictFail   ), //o
    .io_muluIQ_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_exceptionInfo_exception    ), //o
    .io_muluIQ_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_exceptionInfo_eCode[5:0]   ), //o
    .io_muluIQ_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_exceptionInfo_eSubCode     ), //o
    .io_muluIQ_payload_pc                        (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_pc[31:0]                   ), //o
    .io_muluIQ_payload_prd                       (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_prd[5:0]                   ), //o
    .io_muluIQ_payload_psrc_0                    (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_psrc_0[5:0]                ), //o
    .io_muluIQ_payload_psrc_1                    (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_psrc_1[5:0]                ), //o
    .io_muluIQ_payload_imm                       (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_imm[31:0]                  ), //o
    .io_muluIQ_payload_uop_muluOp                (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_uop_muluOp[1:0]            ), //o
    .io_muluIQ_payload_srcReady_0                (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_srcReady_0                 ), //o
    .io_muluIQ_payload_srcReady_1                (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_srcReady_1                 ), //o
    .io_divuIQ_valid                             (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_valid                              ), //o
    .io_divuIQ_ready                             (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_input_ready                           ), //i
    .io_divuIQ_payload_robIdx                    (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_robIdx[4:0]                ), //o
    .io_divuIQ_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_branchResult_targetPC[31:0]), //o
    .io_divuIQ_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_branchResult_branchResult  ), //o
    .io_divuIQ_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_branchResult_predictFail   ), //o
    .io_divuIQ_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_exceptionInfo_exception    ), //o
    .io_divuIQ_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_exceptionInfo_eCode[5:0]   ), //o
    .io_divuIQ_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_exceptionInfo_eSubCode     ), //o
    .io_divuIQ_payload_pc                        (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_pc[31:0]                   ), //o
    .io_divuIQ_payload_prd                       (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_prd[5:0]                   ), //o
    .io_divuIQ_payload_psrc_0                    (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_psrc_0[5:0]                ), //o
    .io_divuIQ_payload_psrc_1                    (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_psrc_1[5:0]                ), //o
    .io_divuIQ_payload_imm                       (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_imm[31:0]                  ), //o
    .io_divuIQ_payload_uop_divuOp                (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_uop_divuOp[1:0]            ), //o
    .io_divuIQ_payload_srcReady_0                (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_srcReady_0                 ), //o
    .io_divuIQ_payload_srcReady_1                (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_srcReady_1                 ), //o
    .io_lsuIQ_valid                              (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_valid                               ), //o
    .io_lsuIQ_ready                              (cpuClockingArea_areaFlushReset_issueQueueLSU_io_input_ready                            ), //i
    .io_lsuIQ_payload_robIdx                     (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_robIdx[4:0]                 ), //o
    .io_lsuIQ_payload_branchResult_targetPC      (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_branchResult_targetPC[31:0] ), //o
    .io_lsuIQ_payload_branchResult_branchResult  (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_branchResult_branchResult   ), //o
    .io_lsuIQ_payload_branchResult_predictFail   (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_branchResult_predictFail    ), //o
    .io_lsuIQ_payload_exceptionInfo_exception    (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_exceptionInfo_exception     ), //o
    .io_lsuIQ_payload_exceptionInfo_eCode        (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_exceptionInfo_eCode[5:0]    ), //o
    .io_lsuIQ_payload_exceptionInfo_eSubCode     (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_exceptionInfo_eSubCode      ), //o
    .io_lsuIQ_payload_pc                         (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_pc[31:0]                    ), //o
    .io_lsuIQ_payload_prd                        (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_prd[5:0]                    ), //o
    .io_lsuIQ_payload_psrc_0                     (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_psrc_0[5:0]                 ), //o
    .io_lsuIQ_payload_psrc_1                     (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_psrc_1[5:0]                 ), //o
    .io_lsuIQ_payload_imm                        (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_imm[31:0]                   ), //o
    .io_lsuIQ_payload_uop_lsuOp                  (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_uop_lsuOp[3:0]              ), //o
    .io_lsuIQ_payload_uop_lsuCoOp                (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_uop_lsuCoOp[4:0]            ), //o
    .io_lsuIQ_payload_roop_lsuROOp               (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_roop_lsuROOp                ), //o
    .io_lsuIQ_payload_srcReady_0                 (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_srcReady_0                  ), //o
    .io_lsuIQ_payload_srcReady_1                 (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_srcReady_1                  )  //o
  );
  IssueQueue cpuClockingArea_areaFlushReset_issueQueueALU0 (
    .io_input_valid                             (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_valid                                 ), //i
    .io_input_ready                             (cpuClockingArea_areaFlushReset_issueQueueALU0_io_input_ready                              ), //o
    .io_input_payload_robIdx                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_robIdx[4:0]                   ), //i
    .io_input_payload_branchInfo_predictPC      (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_branchInfo_predictPC[31:0]    ), //i
    .io_input_payload_branchInfo_predictResult  (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_branchInfo_predictResult      ), //i
    .io_input_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_exceptionInfo_exception       ), //i
    .io_input_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_exceptionInfo_eCode[5:0]      ), //i
    .io_input_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_exceptionInfo_eSubCode        ), //i
    .io_input_payload_pc                        (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_pc[31:0]                      ), //i
    .io_input_payload_prd                       (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_prd[5:0]                      ), //i
    .io_input_payload_psrc_0                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_psrc_0[5:0]                   ), //i
    .io_input_payload_psrc_1                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_psrc_1[5:0]                   ), //i
    .io_input_payload_imm                       (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_imm[31:0]                     ), //i
    .io_input_payload_uop_aluOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_uop_aluOp[3:0]                ), //i
    .io_input_payload_uop_bruOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_uop_bruOp[1:0]                ), //i
    .io_input_payload_uop_cruOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_uop_cruOp[1:0]                ), //i
    .io_input_payload_roop_aluROOp              (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_roop_aluROOp[2:0]             ), //i
    .io_input_payload_srcReady_0                (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_srcReady_0                    ), //i
    .io_input_payload_srcReady_1                (cpuClockingArea_areaFlushReset_dispatcher_io_alu0IQ_payload_srcReady_1                    ), //i
    .io_csrInQueue                              (cpuClockingArea_areaFlushReset_issueQueueALU0_io_csrInQueue                               ), //o
    .io_output_valid                            (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_valid                             ), //o
    .io_output_ready                            (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_ready                             ), //i
    .io_output_payload_robIdx                   (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_robIdx[4:0]               ), //o
    .io_output_payload_branchInfo_predictPC     (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_branchInfo_predictPC[31:0]), //o
    .io_output_payload_branchInfo_predictResult (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_branchInfo_predictResult  ), //o
    .io_output_payload_exceptionInfo_exception  (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_exceptionInfo_exception   ), //o
    .io_output_payload_exceptionInfo_eCode      (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_exceptionInfo_eCode[5:0]  ), //o
    .io_output_payload_exceptionInfo_eSubCode   (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_exceptionInfo_eSubCode    ), //o
    .io_output_payload_pc                       (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_pc[31:0]                  ), //o
    .io_output_payload_prd                      (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_prd[5:0]                  ), //o
    .io_output_payload_psrc_0                   (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_psrc_0[5:0]               ), //o
    .io_output_payload_psrc_1                   (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_psrc_1[5:0]               ), //o
    .io_output_payload_imm                      (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_imm[31:0]                 ), //o
    .io_output_payload_uop_aluOp                (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_uop_aluOp[3:0]            ), //o
    .io_output_payload_uop_bruOp                (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_uop_bruOp[1:0]            ), //o
    .io_output_payload_uop_cruOp                (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_uop_cruOp[1:0]            ), //o
    .io_output_payload_roop_aluROOp             (cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_roop_aluROOp[2:0]         ), //o
    .io_writebackSignal_0                       (cpuClockingArea_areaFlushReset_commitALU0_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_1                       (cpuClockingArea_areaFlushReset_commitALU1_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_2                       (cpuClockingArea_areaFlushReset_commitMULU_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_3                       (cpuClockingArea_areaFlushReset_commitDIVU_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_4                       (cpuClockingArea_areaFlushReset_commitLSU_io_prf_idx[5:0]                                  ), //i
    .io_earlyWakeup_0_valid                     (cpuClockingArea_areaFlushReset_issueQueueALU0_io_wakeOut_valid                            ), //i
    .io_earlyWakeup_0_payload                   (cpuClockingArea_areaFlushReset_issueQueueALU0_io_wakeOut_payload[5:0]                     ), //i
    .io_earlyWakeup_1_valid                     (cpuClockingArea_areaFlushReset_roALU0_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_1_payload                   (cpuClockingArea_areaFlushReset_roALU0_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_2_valid                     (cpuClockingArea_areaFlushReset_fuALU0_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_2_payload                   (cpuClockingArea_areaFlushReset_fuALU0_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_3_valid                     (cpuClockingArea_areaFlushReset_issueQueueALU1_io_wakeOut_valid                            ), //i
    .io_earlyWakeup_3_payload                   (cpuClockingArea_areaFlushReset_issueQueueALU1_io_wakeOut_payload[5:0]                     ), //i
    .io_earlyWakeup_4_valid                     (cpuClockingArea_areaFlushReset_roALU1_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_4_payload                   (cpuClockingArea_areaFlushReset_roALU1_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_5_valid                     (cpuClockingArea_areaFlushReset_fuALU1_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_5_payload                   (cpuClockingArea_areaFlushReset_fuALU1_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_6_valid                     (cpuClockingArea_fuLSU_io_wakeOut_0_valid                                                  ), //i
    .io_earlyWakeup_6_payload                   (cpuClockingArea_fuLSU_io_wakeOut_0_payload[5:0]                                           ), //i
    .io_earlyWakeup_7_valid                     (cpuClockingArea_fuLSU_io_wakeOut_1_valid                                                  ), //i
    .io_earlyWakeup_7_payload                   (cpuClockingArea_fuLSU_io_wakeOut_1_payload[5:0]                                           ), //i
    .io_wakeOut_valid                           (cpuClockingArea_areaFlushReset_issueQueueALU0_io_wakeOut_valid                            ), //o
    .io_wakeOut_payload                         (cpuClockingArea_areaFlushReset_issueQueueALU0_io_wakeOut_payload[5:0]                     ), //o
    .aclk                                       (aclk                                                                                      ), //i
    .cpuClockingArea_areaFlushReset_newReset    (cpuClockingArea_areaFlushReset_newReset                                                   )  //i
  );
  IssueQueue_1 cpuClockingArea_areaFlushReset_issueQueueALU1 (
    .io_input_valid                             (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_valid                                 ), //i
    .io_input_ready                             (cpuClockingArea_areaFlushReset_issueQueueALU1_io_input_ready                              ), //o
    .io_input_payload_robIdx                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_robIdx[4:0]                   ), //i
    .io_input_payload_branchInfo_predictPC      (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_branchInfo_predictPC[31:0]    ), //i
    .io_input_payload_branchInfo_predictResult  (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_branchInfo_predictResult      ), //i
    .io_input_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_exceptionInfo_exception       ), //i
    .io_input_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_exceptionInfo_eCode[5:0]      ), //i
    .io_input_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_exceptionInfo_eSubCode        ), //i
    .io_input_payload_pc                        (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_pc[31:0]                      ), //i
    .io_input_payload_prd                       (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_prd[5:0]                      ), //i
    .io_input_payload_psrc_0                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_psrc_0[5:0]                   ), //i
    .io_input_payload_psrc_1                    (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_psrc_1[5:0]                   ), //i
    .io_input_payload_imm                       (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_imm[31:0]                     ), //i
    .io_input_payload_uop_aluOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_uop_aluOp[3:0]                ), //i
    .io_input_payload_uop_bruOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_uop_bruOp[1:0]                ), //i
    .io_input_payload_roop_aluROOp              (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_roop_aluROOp[2:0]             ), //i
    .io_input_payload_roop_cruROOp              (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_roop_cruROOp[1:0]             ), //i
    .io_input_payload_srcReady_0                (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_srcReady_0                    ), //i
    .io_input_payload_srcReady_1                (cpuClockingArea_areaFlushReset_dispatcher_io_alu1IQ_payload_srcReady_1                    ), //i
    .io_csrInQueue                              (cpuClockingArea_areaFlushReset_issueQueueALU1_io_csrInQueue                               ), //o
    .io_output_valid                            (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_valid                             ), //o
    .io_output_ready                            (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_ready                             ), //i
    .io_output_payload_robIdx                   (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_robIdx[4:0]               ), //o
    .io_output_payload_branchInfo_predictPC     (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_branchInfo_predictPC[31:0]), //o
    .io_output_payload_branchInfo_predictResult (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_branchInfo_predictResult  ), //o
    .io_output_payload_exceptionInfo_exception  (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_exceptionInfo_exception   ), //o
    .io_output_payload_exceptionInfo_eCode      (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_exceptionInfo_eCode[5:0]  ), //o
    .io_output_payload_exceptionInfo_eSubCode   (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_exceptionInfo_eSubCode    ), //o
    .io_output_payload_pc                       (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_pc[31:0]                  ), //o
    .io_output_payload_prd                      (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_prd[5:0]                  ), //o
    .io_output_payload_psrc_0                   (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_psrc_0[5:0]               ), //o
    .io_output_payload_psrc_1                   (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_psrc_1[5:0]               ), //o
    .io_output_payload_imm                      (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_imm[31:0]                 ), //o
    .io_output_payload_uop_aluOp                (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_uop_aluOp[3:0]            ), //o
    .io_output_payload_uop_bruOp                (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_uop_bruOp[1:0]            ), //o
    .io_output_payload_roop_aluROOp             (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_roop_aluROOp[2:0]         ), //o
    .io_output_payload_roop_cruROOp             (cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_roop_cruROOp[1:0]         ), //o
    .io_writebackSignal_0                       (cpuClockingArea_areaFlushReset_commitALU0_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_1                       (cpuClockingArea_areaFlushReset_commitALU1_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_2                       (cpuClockingArea_areaFlushReset_commitMULU_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_3                       (cpuClockingArea_areaFlushReset_commitDIVU_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_4                       (cpuClockingArea_areaFlushReset_commitLSU_io_prf_idx[5:0]                                  ), //i
    .io_earlyWakeup_0_valid                     (cpuClockingArea_areaFlushReset_issueQueueALU0_io_wakeOut_valid                            ), //i
    .io_earlyWakeup_0_payload                   (cpuClockingArea_areaFlushReset_issueQueueALU0_io_wakeOut_payload[5:0]                     ), //i
    .io_earlyWakeup_1_valid                     (cpuClockingArea_areaFlushReset_roALU0_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_1_payload                   (cpuClockingArea_areaFlushReset_roALU0_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_2_valid                     (cpuClockingArea_areaFlushReset_fuALU0_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_2_payload                   (cpuClockingArea_areaFlushReset_fuALU0_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_3_valid                     (cpuClockingArea_areaFlushReset_issueQueueALU1_io_wakeOut_valid                            ), //i
    .io_earlyWakeup_3_payload                   (cpuClockingArea_areaFlushReset_issueQueueALU1_io_wakeOut_payload[5:0]                     ), //i
    .io_earlyWakeup_4_valid                     (cpuClockingArea_areaFlushReset_roALU1_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_4_payload                   (cpuClockingArea_areaFlushReset_roALU1_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_5_valid                     (cpuClockingArea_areaFlushReset_fuALU1_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_5_payload                   (cpuClockingArea_areaFlushReset_fuALU1_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_6_valid                     (cpuClockingArea_fuLSU_io_wakeOut_0_valid                                                  ), //i
    .io_earlyWakeup_6_payload                   (cpuClockingArea_fuLSU_io_wakeOut_0_payload[5:0]                                           ), //i
    .io_earlyWakeup_7_valid                     (cpuClockingArea_fuLSU_io_wakeOut_1_valid                                                  ), //i
    .io_earlyWakeup_7_payload                   (cpuClockingArea_fuLSU_io_wakeOut_1_payload[5:0]                                           ), //i
    .io_wakeOut_valid                           (cpuClockingArea_areaFlushReset_issueQueueALU1_io_wakeOut_valid                            ), //o
    .io_wakeOut_payload                         (cpuClockingArea_areaFlushReset_issueQueueALU1_io_wakeOut_payload[5:0]                     ), //o
    .aclk                                       (aclk                                                                                      ), //i
    .cpuClockingArea_areaFlushReset_newReset    (cpuClockingArea_areaFlushReset_newReset                                                   )  //i
  );
  IssueQueue_2 cpuClockingArea_areaFlushReset_issueQueueMULU (
    .io_input_valid                              (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_valid                                  ), //i
    .io_input_ready                              (cpuClockingArea_areaFlushReset_issueQueueMULU_io_input_ready                               ), //o
    .io_input_payload_robIdx                     (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_robIdx[4:0]                    ), //i
    .io_input_payload_branchResult_targetPC      (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_branchResult_targetPC[31:0]    ), //i
    .io_input_payload_branchResult_branchResult  (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_branchResult_branchResult      ), //i
    .io_input_payload_branchResult_predictFail   (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_branchResult_predictFail       ), //i
    .io_input_payload_exceptionInfo_exception    (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_exceptionInfo_exception        ), //i
    .io_input_payload_exceptionInfo_eCode        (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_exceptionInfo_eCode[5:0]       ), //i
    .io_input_payload_exceptionInfo_eSubCode     (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_exceptionInfo_eSubCode         ), //i
    .io_input_payload_pc                         (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_pc[31:0]                       ), //i
    .io_input_payload_prd                        (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_prd[5:0]                       ), //i
    .io_input_payload_psrc_0                     (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_psrc_0[5:0]                    ), //i
    .io_input_payload_psrc_1                     (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_psrc_1[5:0]                    ), //i
    .io_input_payload_imm                        (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_imm[31:0]                      ), //i
    .io_input_payload_uop_muluOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_uop_muluOp[1:0]                ), //i
    .io_input_payload_srcReady_0                 (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_srcReady_0                     ), //i
    .io_input_payload_srcReady_1                 (cpuClockingArea_areaFlushReset_dispatcher_io_muluIQ_payload_srcReady_1                     ), //i
    .io_output_valid                             (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_valid                              ), //o
    .io_output_ready                             (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_ready                              ), //i
    .io_output_payload_robIdx                    (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_robIdx[4:0]                ), //o
    .io_output_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_branchResult_targetPC[31:0]), //o
    .io_output_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_branchResult_branchResult  ), //o
    .io_output_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_branchResult_predictFail   ), //o
    .io_output_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_exceptionInfo_exception    ), //o
    .io_output_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_exceptionInfo_eCode[5:0]   ), //o
    .io_output_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_exceptionInfo_eSubCode     ), //o
    .io_output_payload_pc                        (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_pc[31:0]                   ), //o
    .io_output_payload_prd                       (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_prd[5:0]                   ), //o
    .io_output_payload_psrc_0                    (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_psrc_0[5:0]                ), //o
    .io_output_payload_psrc_1                    (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_psrc_1[5:0]                ), //o
    .io_output_payload_imm                       (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_imm[31:0]                  ), //o
    .io_output_payload_uop_muluOp                (cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_uop_muluOp[1:0]            ), //o
    .io_writebackSignal_0                        (cpuClockingArea_areaFlushReset_commitALU0_io_prf_idx[5:0]                                  ), //i
    .io_writebackSignal_1                        (cpuClockingArea_areaFlushReset_commitALU1_io_prf_idx[5:0]                                  ), //i
    .io_writebackSignal_2                        (cpuClockingArea_areaFlushReset_commitMULU_io_prf_idx[5:0]                                  ), //i
    .io_writebackSignal_3                        (cpuClockingArea_areaFlushReset_commitDIVU_io_prf_idx[5:0]                                  ), //i
    .io_writebackSignal_4                        (cpuClockingArea_areaFlushReset_commitLSU_io_prf_idx[5:0]                                   ), //i
    .io_earlyWakeup_0_valid                      (cpuClockingArea_fuLSU_io_wakeOut_0_valid                                                   ), //i
    .io_earlyWakeup_0_payload                    (cpuClockingArea_fuLSU_io_wakeOut_0_payload[5:0]                                            ), //i
    .io_earlyWakeup_1_valid                      (cpuClockingArea_fuLSU_io_wakeOut_1_valid                                                   ), //i
    .io_earlyWakeup_1_payload                    (cpuClockingArea_fuLSU_io_wakeOut_1_payload[5:0]                                            ), //i
    .aclk                                        (aclk                                                                                       ), //i
    .cpuClockingArea_areaFlushReset_newReset     (cpuClockingArea_areaFlushReset_newReset                                                    )  //i
  );
  IssueQueue_3 cpuClockingArea_areaFlushReset_issueQueueDIVU (
    .io_input_valid                              (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_valid                                  ), //i
    .io_input_ready                              (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_input_ready                               ), //o
    .io_input_payload_robIdx                     (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_robIdx[4:0]                    ), //i
    .io_input_payload_branchResult_targetPC      (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_branchResult_targetPC[31:0]    ), //i
    .io_input_payload_branchResult_branchResult  (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_branchResult_branchResult      ), //i
    .io_input_payload_branchResult_predictFail   (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_branchResult_predictFail       ), //i
    .io_input_payload_exceptionInfo_exception    (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_exceptionInfo_exception        ), //i
    .io_input_payload_exceptionInfo_eCode        (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_exceptionInfo_eCode[5:0]       ), //i
    .io_input_payload_exceptionInfo_eSubCode     (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_exceptionInfo_eSubCode         ), //i
    .io_input_payload_pc                         (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_pc[31:0]                       ), //i
    .io_input_payload_prd                        (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_prd[5:0]                       ), //i
    .io_input_payload_psrc_0                     (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_psrc_0[5:0]                    ), //i
    .io_input_payload_psrc_1                     (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_psrc_1[5:0]                    ), //i
    .io_input_payload_imm                        (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_imm[31:0]                      ), //i
    .io_input_payload_uop_divuOp                 (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_uop_divuOp[1:0]                ), //i
    .io_input_payload_srcReady_0                 (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_srcReady_0                     ), //i
    .io_input_payload_srcReady_1                 (cpuClockingArea_areaFlushReset_dispatcher_io_divuIQ_payload_srcReady_1                     ), //i
    .io_output_valid                             (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_valid                              ), //o
    .io_output_ready                             (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_ready                              ), //i
    .io_output_payload_robIdx                    (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_robIdx[4:0]                ), //o
    .io_output_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_branchResult_targetPC[31:0]), //o
    .io_output_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_branchResult_branchResult  ), //o
    .io_output_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_branchResult_predictFail   ), //o
    .io_output_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_exceptionInfo_exception    ), //o
    .io_output_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_exceptionInfo_eCode[5:0]   ), //o
    .io_output_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_exceptionInfo_eSubCode     ), //o
    .io_output_payload_pc                        (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_pc[31:0]                   ), //o
    .io_output_payload_prd                       (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_prd[5:0]                   ), //o
    .io_output_payload_psrc_0                    (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_psrc_0[5:0]                ), //o
    .io_output_payload_psrc_1                    (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_psrc_1[5:0]                ), //o
    .io_output_payload_imm                       (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_imm[31:0]                  ), //o
    .io_output_payload_uop_divuOp                (cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_uop_divuOp[1:0]            ), //o
    .io_writebackSignal_0                        (cpuClockingArea_areaFlushReset_commitALU0_io_prf_idx[5:0]                                  ), //i
    .io_writebackSignal_1                        (cpuClockingArea_areaFlushReset_commitALU1_io_prf_idx[5:0]                                  ), //i
    .io_writebackSignal_2                        (cpuClockingArea_areaFlushReset_commitMULU_io_prf_idx[5:0]                                  ), //i
    .io_writebackSignal_3                        (cpuClockingArea_areaFlushReset_commitDIVU_io_prf_idx[5:0]                                  ), //i
    .io_writebackSignal_4                        (cpuClockingArea_areaFlushReset_commitLSU_io_prf_idx[5:0]                                   ), //i
    .aclk                                        (aclk                                                                                       ), //i
    .cpuClockingArea_areaFlushReset_newReset     (cpuClockingArea_areaFlushReset_newReset                                                    )  //i
  );
  IssueQueue_4 cpuClockingArea_areaFlushReset_issueQueueLSU (
    .io_input_valid                              (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_valid                                  ), //i
    .io_input_ready                              (cpuClockingArea_areaFlushReset_issueQueueLSU_io_input_ready                               ), //o
    .io_input_payload_robIdx                     (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_robIdx[4:0]                    ), //i
    .io_input_payload_branchResult_targetPC      (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_branchResult_targetPC[31:0]    ), //i
    .io_input_payload_branchResult_branchResult  (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_branchResult_branchResult      ), //i
    .io_input_payload_branchResult_predictFail   (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_branchResult_predictFail       ), //i
    .io_input_payload_exceptionInfo_exception    (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_exceptionInfo_exception        ), //i
    .io_input_payload_exceptionInfo_eCode        (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_exceptionInfo_eCode[5:0]       ), //i
    .io_input_payload_exceptionInfo_eSubCode     (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_exceptionInfo_eSubCode         ), //i
    .io_input_payload_pc                         (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_pc[31:0]                       ), //i
    .io_input_payload_prd                        (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_prd[5:0]                       ), //i
    .io_input_payload_psrc_0                     (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_psrc_0[5:0]                    ), //i
    .io_input_payload_psrc_1                     (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_psrc_1[5:0]                    ), //i
    .io_input_payload_imm                        (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_imm[31:0]                      ), //i
    .io_input_payload_uop_lsuOp                  (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_uop_lsuOp[3:0]                 ), //i
    .io_input_payload_uop_lsuCoOp                (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_uop_lsuCoOp[4:0]               ), //i
    .io_input_payload_roop_lsuROOp               (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_roop_lsuROOp                   ), //i
    .io_input_payload_srcReady_0                 (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_srcReady_0                     ), //i
    .io_input_payload_srcReady_1                 (cpuClockingArea_areaFlushReset_dispatcher_io_lsuIQ_payload_srcReady_1                     ), //i
    .io_output_valid                             (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_valid                              ), //o
    .io_output_ready                             (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_ready                              ), //i
    .io_output_payload_robIdx                    (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_robIdx[4:0]                ), //o
    .io_output_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_branchResult_targetPC[31:0]), //o
    .io_output_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_branchResult_branchResult  ), //o
    .io_output_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_branchResult_predictFail   ), //o
    .io_output_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_exceptionInfo_exception    ), //o
    .io_output_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_exceptionInfo_eCode[5:0]   ), //o
    .io_output_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_exceptionInfo_eSubCode     ), //o
    .io_output_payload_pc                        (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_pc[31:0]                   ), //o
    .io_output_payload_prd                       (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_prd[5:0]                   ), //o
    .io_output_payload_psrc_0                    (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_psrc_0[5:0]                ), //o
    .io_output_payload_psrc_1                    (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_psrc_1[5:0]                ), //o
    .io_output_payload_imm                       (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_imm[31:0]                  ), //o
    .io_output_payload_uop_lsuOp                 (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_uop_lsuOp[3:0]             ), //o
    .io_output_payload_uop_lsuCoOp               (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_uop_lsuCoOp[4:0]           ), //o
    .io_output_payload_roop_lsuROOp              (cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_roop_lsuROOp               ), //o
    .io_writebackSignal_0                        (cpuClockingArea_areaFlushReset_commitALU0_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_1                        (cpuClockingArea_areaFlushReset_commitALU1_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_2                        (cpuClockingArea_areaFlushReset_commitMULU_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_3                        (cpuClockingArea_areaFlushReset_commitDIVU_io_prf_idx[5:0]                                 ), //i
    .io_writebackSignal_4                        (cpuClockingArea_areaFlushReset_commitLSU_io_prf_idx[5:0]                                  ), //i
    .io_earlyWakeup_0_valid                      (cpuClockingArea_areaFlushReset_issueQueueALU0_io_wakeOut_valid                            ), //i
    .io_earlyWakeup_0_payload                    (cpuClockingArea_areaFlushReset_issueQueueALU0_io_wakeOut_payload[5:0]                     ), //i
    .io_earlyWakeup_1_valid                      (cpuClockingArea_areaFlushReset_roALU0_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_1_payload                    (cpuClockingArea_areaFlushReset_roALU0_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_2_valid                      (cpuClockingArea_areaFlushReset_fuALU0_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_2_payload                    (cpuClockingArea_areaFlushReset_fuALU0_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_3_valid                      (cpuClockingArea_areaFlushReset_issueQueueALU1_io_wakeOut_valid                            ), //i
    .io_earlyWakeup_3_payload                    (cpuClockingArea_areaFlushReset_issueQueueALU1_io_wakeOut_payload[5:0]                     ), //i
    .io_earlyWakeup_4_valid                      (cpuClockingArea_areaFlushReset_roALU1_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_4_payload                    (cpuClockingArea_areaFlushReset_roALU1_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_5_valid                      (cpuClockingArea_areaFlushReset_fuALU1_io_wakeOut_valid                                    ), //i
    .io_earlyWakeup_5_payload                    (cpuClockingArea_areaFlushReset_fuALU1_io_wakeOut_payload[5:0]                             ), //i
    .io_earlyWakeup_6_valid                      (cpuClockingArea_fuLSU_io_wakeOut_0_valid                                                  ), //i
    .io_earlyWakeup_6_payload                    (cpuClockingArea_fuLSU_io_wakeOut_0_payload[5:0]                                           ), //i
    .io_earlyWakeup_7_valid                      (cpuClockingArea_fuLSU_io_wakeOut_1_valid                                                  ), //i
    .io_earlyWakeup_7_payload                    (cpuClockingArea_fuLSU_io_wakeOut_1_payload[5:0]                                           ), //i
    .io_earlyWakeup_8_valid                      (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_0_valid                                  ), //i
    .io_earlyWakeup_8_payload                    (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_0_payload[5:0]                           ), //i
    .io_earlyWakeup_9_valid                      (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_1_valid                                  ), //i
    .io_earlyWakeup_9_payload                    (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_1_payload[5:0]                           ), //i
    .io_earlyWakeup_10_valid                     (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_2_valid                                  ), //i
    .io_earlyWakeup_10_payload                   (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_2_payload[5:0]                           ), //i
    .aclk                                        (aclk                                                                                      ), //i
    .cpuClockingArea_areaFlushReset_newReset     (cpuClockingArea_areaFlushReset_newReset                                                   )  //i
  );
  ReadOperandLogic cpuClockingArea_areaFlushReset_roALU0 (
    .io_cmd_valid                             (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_valid                             ), //i
    .io_cmd_ready                             (cpuClockingArea_areaFlushReset_roALU0_io_cmd_ready                                                         ), //o
    .io_cmd_payload_robIdx                    (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_robIdx[4:0]               ), //i
    .io_cmd_payload_branchInfo_predictPC      (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_branchInfo_predictPC[31:0]), //i
    .io_cmd_payload_branchInfo_predictResult  (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_branchInfo_predictResult  ), //i
    .io_cmd_payload_exceptionInfo_exception   (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_exceptionInfo_exception   ), //i
    .io_cmd_payload_exceptionInfo_eCode       (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_exceptionInfo_eCode[5:0]  ), //i
    .io_cmd_payload_exceptionInfo_eSubCode    (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_exceptionInfo_eSubCode    ), //i
    .io_cmd_payload_pc                        (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_pc[31:0]                  ), //i
    .io_cmd_payload_prd                       (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_prd[5:0]                  ), //i
    .io_cmd_payload_psrc_0                    (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_psrc_0[5:0]               ), //i
    .io_cmd_payload_psrc_1                    (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_psrc_1[5:0]               ), //i
    .io_cmd_payload_imm                       (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_imm[31:0]                 ), //i
    .io_cmd_payload_uop_aluOp                 (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp[3:0]            ), //i
    .io_cmd_payload_uop_bruOp                 (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_bruOp[1:0]            ), //i
    .io_cmd_payload_uop_cruOp                 (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_cruOp[1:0]            ), //i
    .io_cmd_payload_roop_aluROOp              (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp[2:0]         ), //i
    .io_toFU_valid                            (cpuClockingArea_areaFlushReset_roALU0_io_toFU_valid                                                        ), //o
    .io_toFU_ready                            (cpuClockingArea_areaFlushReset_roALU0_io_toFU_ready                                                        ), //i
    .io_toFU_payload_src1                     (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src1[31:0]                                           ), //o
    .io_toFU_payload_src2                     (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src2[31:0]                                           ), //o
    .io_toFU_payload_src3                     (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src3[31:0]                                           ), //o
    .io_toFU_payload_src4                     (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src4[31:0]                                           ), //o
    .io_toFU_payload_robIdx                   (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_robIdx[4:0]                                          ), //o
    .io_toFU_payload_branchInfo_predictPC     (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_branchInfo_predictPC[31:0]                           ), //o
    .io_toFU_payload_branchInfo_predictResult (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_branchInfo_predictResult                             ), //o
    .io_toFU_payload_exceptionInfo_exception  (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_exceptionInfo_exception                              ), //o
    .io_toFU_payload_exceptionInfo_eCode      (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_exceptionInfo_eCode[5:0]                             ), //o
    .io_toFU_payload_exceptionInfo_eSubCode   (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_exceptionInfo_eSubCode                               ), //o
    .io_toFU_payload_pc                       (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_pc[31:0]                                             ), //o
    .io_toFU_payload_prd                      (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_prd[5:0]                                             ), //o
    .io_toFU_payload_uop_aluOp                (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_uop_aluOp[3:0]                                       ), //o
    .io_toFU_payload_uop_bruOp                (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_uop_bruOp[1:0]                                       ), //o
    .io_toFU_payload_uop_cruOp                (cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_uop_cruOp[1:0]                                       ), //o
    .io_forward_0_valid                       (cpuClockingArea_areaFlushReset_fuALU0_io_forward_valid                                                     ), //i
    .io_forward_0_payload_idx                 (cpuClockingArea_areaFlushReset_fuALU0_io_forward_payload_idx[5:0]                                          ), //i
    .io_forward_0_payload_payload             (cpuClockingArea_areaFlushReset_fuALU0_io_forward_payload_payload[31:0]                                     ), //i
    .io_forward_1_valid                       (cpuClockingArea_areaFlushReset_commitALU0_io_forward_valid                                                 ), //i
    .io_forward_1_payload_idx                 (cpuClockingArea_areaFlushReset_commitALU0_io_forward_payload_idx[5:0]                                      ), //i
    .io_forward_1_payload_payload             (cpuClockingArea_areaFlushReset_commitALU0_io_forward_payload_payload[31:0]                                 ), //i
    .io_forward_2_valid                       (cpuClockingArea_areaFlushReset_fuALU1_io_forward_valid                                                     ), //i
    .io_forward_2_payload_idx                 (cpuClockingArea_areaFlushReset_fuALU1_io_forward_payload_idx[5:0]                                          ), //i
    .io_forward_2_payload_payload             (cpuClockingArea_areaFlushReset_fuALU1_io_forward_payload_payload[31:0]                                     ), //i
    .io_forward_3_valid                       (cpuClockingArea_areaFlushReset_commitALU1_io_forward_valid                                                 ), //i
    .io_forward_3_payload_idx                 (cpuClockingArea_areaFlushReset_commitALU1_io_forward_payload_idx[5:0]                                      ), //i
    .io_forward_3_payload_payload             (cpuClockingArea_areaFlushReset_commitALU1_io_forward_payload_payload[31:0]                                 ), //i
    .io_forward_4_valid                       (cpuClockingArea_areaFlushReset_commitLSU_io_forward_valid                                                  ), //i
    .io_forward_4_payload_idx                 (cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_idx[5:0]                                       ), //i
    .io_forward_4_payload_payload             (cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_payload[31:0]                                  ), //i
    .io_wakeOut_valid                         (cpuClockingArea_areaFlushReset_roALU0_io_wakeOut_valid                                                     ), //o
    .io_wakeOut_payload                       (cpuClockingArea_areaFlushReset_roALU0_io_wakeOut_payload[5:0]                                              ), //o
    .io_prf_0_idx                             (cpuClockingArea_areaFlushReset_roALU0_io_prf_0_idx[5:0]                                                    ), //o
    .io_prf_0_data                            (cpuClockingArea_prf_io_read_0_0_data[31:0]                                                                 ), //i
    .io_prf_1_idx                             (cpuClockingArea_areaFlushReset_roALU0_io_prf_1_idx[5:0]                                                    ), //o
    .io_prf_1_data                            (cpuClockingArea_prf_io_read_0_1_data[31:0]                                                                 ), //i
    .io_csr_value                             (cpuClockingArea_csr_io_swRead_value[31:0]                                                                  ), //i
    .io_csr_address                           (cpuClockingArea_areaFlushReset_roALU0_io_csr_address[13:0]                                                 ), //o
    .io_interrupt                             (cpuClockingArea_csr_io_interrupt                                                                           )  //i
  );
  ReadOperandLogic_1 cpuClockingArea_areaFlushReset_roALU1 (
    .io_cmd_valid                             (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_valid                             ), //i
    .io_cmd_ready                             (cpuClockingArea_areaFlushReset_roALU1_io_cmd_ready                                                         ), //o
    .io_cmd_payload_robIdx                    (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_robIdx[4:0]               ), //i
    .io_cmd_payload_branchInfo_predictPC      (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_branchInfo_predictPC[31:0]), //i
    .io_cmd_payload_branchInfo_predictResult  (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_branchInfo_predictResult  ), //i
    .io_cmd_payload_exceptionInfo_exception   (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_exceptionInfo_exception   ), //i
    .io_cmd_payload_exceptionInfo_eCode       (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_exceptionInfo_eCode[5:0]  ), //i
    .io_cmd_payload_exceptionInfo_eSubCode    (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_exceptionInfo_eSubCode    ), //i
    .io_cmd_payload_pc                        (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_pc[31:0]                  ), //i
    .io_cmd_payload_prd                       (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_prd[5:0]                  ), //i
    .io_cmd_payload_psrc_0                    (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_psrc_0[5:0]               ), //i
    .io_cmd_payload_psrc_1                    (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_psrc_1[5:0]               ), //i
    .io_cmd_payload_imm                       (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_imm[31:0]                 ), //i
    .io_cmd_payload_uop_aluOp                 (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp[3:0]            ), //i
    .io_cmd_payload_uop_bruOp                 (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_bruOp[1:0]            ), //i
    .io_cmd_payload_roop_aluROOp              (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp[2:0]         ), //i
    .io_cmd_payload_roop_cruROOp              (toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_cruROOp[1:0]         ), //i
    .io_toFU_valid                            (cpuClockingArea_areaFlushReset_roALU1_io_toFU_valid                                                        ), //o
    .io_toFU_ready                            (cpuClockingArea_areaFlushReset_roALU1_io_toFU_ready                                                        ), //i
    .io_toFU_payload_src1                     (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src1[31:0]                                           ), //o
    .io_toFU_payload_src2                     (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src2[31:0]                                           ), //o
    .io_toFU_payload_src3                     (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src3[31:0]                                           ), //o
    .io_toFU_payload_src4                     (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src4[31:0]                                           ), //o
    .io_toFU_payload_robIdx                   (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_robIdx[4:0]                                          ), //o
    .io_toFU_payload_branchInfo_predictPC     (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_branchInfo_predictPC[31:0]                           ), //o
    .io_toFU_payload_branchInfo_predictResult (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_branchInfo_predictResult                             ), //o
    .io_toFU_payload_exceptionInfo_exception  (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_exceptionInfo_exception                              ), //o
    .io_toFU_payload_exceptionInfo_eCode      (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_exceptionInfo_eCode[5:0]                             ), //o
    .io_toFU_payload_exceptionInfo_eSubCode   (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_exceptionInfo_eSubCode                               ), //o
    .io_toFU_payload_pc                       (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_pc[31:0]                                             ), //o
    .io_toFU_payload_prd                      (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_prd[5:0]                                             ), //o
    .io_toFU_payload_uop_aluOp                (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_uop_aluOp[3:0]                                       ), //o
    .io_toFU_payload_uop_bruOp                (cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_uop_bruOp[1:0]                                       ), //o
    .io_forward_0_valid                       (cpuClockingArea_areaFlushReset_fuALU0_io_forward_valid                                                     ), //i
    .io_forward_0_payload_idx                 (cpuClockingArea_areaFlushReset_fuALU0_io_forward_payload_idx[5:0]                                          ), //i
    .io_forward_0_payload_payload             (cpuClockingArea_areaFlushReset_fuALU0_io_forward_payload_payload[31:0]                                     ), //i
    .io_forward_1_valid                       (cpuClockingArea_areaFlushReset_commitALU0_io_forward_valid                                                 ), //i
    .io_forward_1_payload_idx                 (cpuClockingArea_areaFlushReset_commitALU0_io_forward_payload_idx[5:0]                                      ), //i
    .io_forward_1_payload_payload             (cpuClockingArea_areaFlushReset_commitALU0_io_forward_payload_payload[31:0]                                 ), //i
    .io_forward_2_valid                       (cpuClockingArea_areaFlushReset_fuALU1_io_forward_valid                                                     ), //i
    .io_forward_2_payload_idx                 (cpuClockingArea_areaFlushReset_fuALU1_io_forward_payload_idx[5:0]                                          ), //i
    .io_forward_2_payload_payload             (cpuClockingArea_areaFlushReset_fuALU1_io_forward_payload_payload[31:0]                                     ), //i
    .io_forward_3_valid                       (cpuClockingArea_areaFlushReset_commitALU1_io_forward_valid                                                 ), //i
    .io_forward_3_payload_idx                 (cpuClockingArea_areaFlushReset_commitALU1_io_forward_payload_idx[5:0]                                      ), //i
    .io_forward_3_payload_payload             (cpuClockingArea_areaFlushReset_commitALU1_io_forward_payload_payload[31:0]                                 ), //i
    .io_forward_4_valid                       (cpuClockingArea_areaFlushReset_commitLSU_io_forward_valid                                                  ), //i
    .io_forward_4_payload_idx                 (cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_idx[5:0]                                       ), //i
    .io_forward_4_payload_payload             (cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_payload[31:0]                                  ), //i
    .io_wakeOut_valid                         (cpuClockingArea_areaFlushReset_roALU1_io_wakeOut_valid                                                     ), //o
    .io_wakeOut_payload                       (cpuClockingArea_areaFlushReset_roALU1_io_wakeOut_payload[5:0]                                              ), //o
    .io_prf_0_idx                             (cpuClockingArea_areaFlushReset_roALU1_io_prf_0_idx[5:0]                                                    ), //o
    .io_prf_0_data                            (cpuClockingArea_prf_io_read_1_0_data[31:0]                                                                 ), //i
    .io_prf_1_idx                             (cpuClockingArea_areaFlushReset_roALU1_io_prf_1_idx[5:0]                                                    ), //o
    .io_prf_1_data                            (cpuClockingArea_prf_io_read_1_1_data[31:0]                                                                 ), //i
    .io_counter_id                            (cpuClockingArea_csr_io_counter_id[31:0]                                                                    ), //i
    .io_counter_value                         (cpuClockingArea_csr_io_counter_value[63:0]                                                                 ), //i
    .io_interrupt                             (cpuClockingArea_csr_io_interrupt                                                                           )  //i
  );
  ReadOperandLogic_2 cpuClockingArea_areaFlushReset_roMULU (
    .io_cmd_valid                              (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_valid                              ), //i
    .io_cmd_ready                              (cpuClockingArea_areaFlushReset_roMULU_io_cmd_ready                                                          ), //o
    .io_cmd_payload_robIdx                     (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_robIdx[4:0]                ), //i
    .io_cmd_payload_branchResult_targetPC      (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_branchResult_targetPC[31:0]), //i
    .io_cmd_payload_branchResult_branchResult  (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_branchResult_branchResult  ), //i
    .io_cmd_payload_branchResult_predictFail   (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_branchResult_predictFail   ), //i
    .io_cmd_payload_exceptionInfo_exception    (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_exceptionInfo_exception    ), //i
    .io_cmd_payload_exceptionInfo_eCode        (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_exceptionInfo_eCode[5:0]   ), //i
    .io_cmd_payload_exceptionInfo_eSubCode     (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_exceptionInfo_eSubCode     ), //i
    .io_cmd_payload_pc                         (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_pc[31:0]                   ), //i
    .io_cmd_payload_prd                        (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_prd[5:0]                   ), //i
    .io_cmd_payload_psrc_0                     (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_psrc_0[5:0]                ), //i
    .io_cmd_payload_psrc_1                     (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_psrc_1[5:0]                ), //i
    .io_cmd_payload_imm                        (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_imm[31:0]                  ), //i
    .io_cmd_payload_uop_muluOp                 (toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_uop_muluOp[1:0]            ), //i
    .io_toFU_valid                             (cpuClockingArea_areaFlushReset_roMULU_io_toFU_valid                                                         ), //o
    .io_toFU_ready                             (cpuClockingArea_areaFlushReset_roMULU_io_toFU_ready                                                         ), //i
    .io_toFU_payload_src1                      (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_src1[31:0]                                            ), //o
    .io_toFU_payload_src2                      (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_src2[31:0]                                            ), //o
    .io_toFU_payload_robIdx                    (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_robIdx[4:0]                                           ), //o
    .io_toFU_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_branchResult_targetPC[31:0]                           ), //o
    .io_toFU_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_branchResult_branchResult                             ), //o
    .io_toFU_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_branchResult_predictFail                              ), //o
    .io_toFU_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_exceptionInfo_exception                               ), //o
    .io_toFU_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_exceptionInfo_eCode[5:0]                              ), //o
    .io_toFU_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_exceptionInfo_eSubCode                                ), //o
    .io_toFU_payload_pc                        (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_pc[31:0]                                              ), //o
    .io_toFU_payload_prd                       (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_prd[5:0]                                              ), //o
    .io_toFU_payload_uop_muluOp                (cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_uop_muluOp[1:0]                                       ), //o
    .io_forward_0_valid                        (cpuClockingArea_areaFlushReset_commitLSU_io_forward_valid                                                   ), //i
    .io_forward_0_payload_idx                  (cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_idx[5:0]                                        ), //i
    .io_forward_0_payload_payload              (cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_payload[31:0]                                   ), //i
    .io_prf_0_idx                              (cpuClockingArea_areaFlushReset_roMULU_io_prf_0_idx[5:0]                                                     ), //o
    .io_prf_0_data                             (cpuClockingArea_prf_io_read_2_0_data[31:0]                                                                  ), //i
    .io_prf_1_idx                              (cpuClockingArea_areaFlushReset_roMULU_io_prf_1_idx[5:0]                                                     ), //o
    .io_prf_1_data                             (cpuClockingArea_prf_io_read_2_1_data[31:0]                                                                  ), //i
    .io_interrupt                              (cpuClockingArea_csr_io_interrupt                                                                            )  //i
  );
  ReadOperandLogic_3 cpuClockingArea_areaFlushReset_roDIVU (
    .io_cmd_valid                              (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_valid                              ), //i
    .io_cmd_ready                              (cpuClockingArea_areaFlushReset_roDIVU_io_cmd_ready                                                          ), //o
    .io_cmd_payload_robIdx                     (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_robIdx[4:0]                ), //i
    .io_cmd_payload_branchResult_targetPC      (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_branchResult_targetPC[31:0]), //i
    .io_cmd_payload_branchResult_branchResult  (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_branchResult_branchResult  ), //i
    .io_cmd_payload_branchResult_predictFail   (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_branchResult_predictFail   ), //i
    .io_cmd_payload_exceptionInfo_exception    (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_exceptionInfo_exception    ), //i
    .io_cmd_payload_exceptionInfo_eCode        (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_exceptionInfo_eCode[5:0]   ), //i
    .io_cmd_payload_exceptionInfo_eSubCode     (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_exceptionInfo_eSubCode     ), //i
    .io_cmd_payload_pc                         (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_pc[31:0]                   ), //i
    .io_cmd_payload_prd                        (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_prd[5:0]                   ), //i
    .io_cmd_payload_psrc_0                     (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_psrc_0[5:0]                ), //i
    .io_cmd_payload_psrc_1                     (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_psrc_1[5:0]                ), //i
    .io_cmd_payload_imm                        (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_imm[31:0]                  ), //i
    .io_cmd_payload_uop_divuOp                 (toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_uop_divuOp[1:0]            ), //i
    .io_toFU_valid                             (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_valid                                                         ), //o
    .io_toFU_ready                             (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_ready                                                         ), //i
    .io_toFU_payload_src1                      (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_src1[31:0]                                            ), //o
    .io_toFU_payload_src2                      (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_src2[31:0]                                            ), //o
    .io_toFU_payload_robIdx                    (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_robIdx[4:0]                                           ), //o
    .io_toFU_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_branchResult_targetPC[31:0]                           ), //o
    .io_toFU_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_branchResult_branchResult                             ), //o
    .io_toFU_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_branchResult_predictFail                              ), //o
    .io_toFU_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_exceptionInfo_exception                               ), //o
    .io_toFU_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_exceptionInfo_eCode[5:0]                              ), //o
    .io_toFU_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_exceptionInfo_eSubCode                                ), //o
    .io_toFU_payload_pc                        (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_pc[31:0]                                              ), //o
    .io_toFU_payload_prd                       (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_prd[5:0]                                              ), //o
    .io_toFU_payload_uop_divuOp                (cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_uop_divuOp[1:0]                                       ), //o
    .io_prf_0_idx                              (cpuClockingArea_areaFlushReset_roDIVU_io_prf_0_idx[5:0]                                                     ), //o
    .io_prf_0_data                             (cpuClockingArea_prf_io_read_3_0_data[31:0]                                                                  ), //i
    .io_prf_1_idx                              (cpuClockingArea_areaFlushReset_roDIVU_io_prf_1_idx[5:0]                                                     ), //o
    .io_prf_1_data                             (cpuClockingArea_prf_io_read_3_1_data[31:0]                                                                  ), //i
    .io_interrupt                              (cpuClockingArea_csr_io_interrupt                                                                            )  //i
  );
  ReadOperandLogic_4 cpuClockingArea_areaFlushReset_roLSU (
    .io_cmd_valid                              (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_valid                              ), //i
    .io_cmd_ready                              (cpuClockingArea_areaFlushReset_roLSU_io_cmd_ready                                                          ), //o
    .io_cmd_payload_robIdx                     (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_robIdx[4:0]                ), //i
    .io_cmd_payload_branchResult_targetPC      (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_branchResult_targetPC[31:0]), //i
    .io_cmd_payload_branchResult_branchResult  (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_branchResult_branchResult  ), //i
    .io_cmd_payload_branchResult_predictFail   (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_branchResult_predictFail   ), //i
    .io_cmd_payload_exceptionInfo_exception    (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_exceptionInfo_exception    ), //i
    .io_cmd_payload_exceptionInfo_eCode        (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_exceptionInfo_eCode[5:0]   ), //i
    .io_cmd_payload_exceptionInfo_eSubCode     (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_exceptionInfo_eSubCode     ), //i
    .io_cmd_payload_pc                         (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_pc[31:0]                   ), //i
    .io_cmd_payload_prd                        (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_prd[5:0]                   ), //i
    .io_cmd_payload_psrc_0                     (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_psrc_0[5:0]                ), //i
    .io_cmd_payload_psrc_1                     (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_psrc_1[5:0]                ), //i
    .io_cmd_payload_imm                        (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_imm[31:0]                  ), //i
    .io_cmd_payload_uop_lsuOp                  (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp[3:0]             ), //i
    .io_cmd_payload_uop_lsuCoOp                (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuCoOp[4:0]           ), //i
    .io_cmd_payload_roop_lsuROOp               (toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_roop_lsuROOp               ), //i
    .io_toFU_valid                             (cpuClockingArea_areaFlushReset_roLSU_io_toFU_valid                                                         ), //o
    .io_toFU_ready                             (cpuClockingArea_areaFlushReset_roLSU_io_toFU_ready                                                         ), //i
    .io_toFU_payload_src1                      (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_src1[31:0]                                            ), //o
    .io_toFU_payload_src2                      (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_src2[31:0]                                            ), //o
    .io_toFU_payload_src3                      (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_src3[31:0]                                            ), //o
    .io_toFU_payload_robIdx                    (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_robIdx[4:0]                                           ), //o
    .io_toFU_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_branchResult_targetPC[31:0]                           ), //o
    .io_toFU_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_branchResult_branchResult                             ), //o
    .io_toFU_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_branchResult_predictFail                              ), //o
    .io_toFU_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_exceptionInfo_exception                               ), //o
    .io_toFU_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_exceptionInfo_eCode[5:0]                              ), //o
    .io_toFU_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_exceptionInfo_eSubCode                                ), //o
    .io_toFU_payload_pc                        (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_pc[31:0]                                              ), //o
    .io_toFU_payload_prd                       (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_prd[5:0]                                              ), //o
    .io_toFU_payload_uop_lsuOp                 (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_uop_lsuOp[3:0]                                        ), //o
    .io_toFU_payload_uop_lsuCoOp               (cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_uop_lsuCoOp[4:0]                                      ), //o
    .io_forward_0_valid                        (cpuClockingArea_areaFlushReset_fuALU0_io_forward_valid                                                     ), //i
    .io_forward_0_payload_idx                  (cpuClockingArea_areaFlushReset_fuALU0_io_forward_payload_idx[5:0]                                          ), //i
    .io_forward_0_payload_payload              (cpuClockingArea_areaFlushReset_fuALU0_io_forward_payload_payload[31:0]                                     ), //i
    .io_forward_1_valid                        (cpuClockingArea_areaFlushReset_commitALU0_io_forward_valid                                                 ), //i
    .io_forward_1_payload_idx                  (cpuClockingArea_areaFlushReset_commitALU0_io_forward_payload_idx[5:0]                                      ), //i
    .io_forward_1_payload_payload              (cpuClockingArea_areaFlushReset_commitALU0_io_forward_payload_payload[31:0]                                 ), //i
    .io_forward_2_valid                        (cpuClockingArea_areaFlushReset_fuALU1_io_forward_valid                                                     ), //i
    .io_forward_2_payload_idx                  (cpuClockingArea_areaFlushReset_fuALU1_io_forward_payload_idx[5:0]                                          ), //i
    .io_forward_2_payload_payload              (cpuClockingArea_areaFlushReset_fuALU1_io_forward_payload_payload[31:0]                                     ), //i
    .io_forward_3_valid                        (cpuClockingArea_areaFlushReset_commitALU1_io_forward_valid                                                 ), //i
    .io_forward_3_payload_idx                  (cpuClockingArea_areaFlushReset_commitALU1_io_forward_payload_idx[5:0]                                      ), //i
    .io_forward_3_payload_payload              (cpuClockingArea_areaFlushReset_commitALU1_io_forward_payload_payload[31:0]                                 ), //i
    .io_forward_4_valid                        (cpuClockingArea_areaFlushReset_commitLSU_io_forward_valid                                                  ), //i
    .io_forward_4_payload_idx                  (cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_idx[5:0]                                       ), //i
    .io_forward_4_payload_payload              (cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_payload[31:0]                                  ), //i
    .io_forward_5_valid                        (cpuClockingArea_areaFlushReset_fuMULU_io_forward_valid                                                     ), //i
    .io_forward_5_payload_idx                  (cpuClockingArea_areaFlushReset_fuMULU_io_forward_payload_idx[5:0]                                          ), //i
    .io_forward_5_payload_payload              (cpuClockingArea_areaFlushReset_fuMULU_io_forward_payload_payload[31:0]                                     ), //i
    .io_forward_6_valid                        (cpuClockingArea_areaFlushReset_commitMULU_io_forward_valid                                                 ), //i
    .io_forward_6_payload_idx                  (cpuClockingArea_areaFlushReset_commitMULU_io_forward_payload_idx[5:0]                                      ), //i
    .io_forward_6_payload_payload              (cpuClockingArea_areaFlushReset_commitMULU_io_forward_payload_payload[31:0]                                 ), //i
    .io_prf_0_idx                              (cpuClockingArea_areaFlushReset_roLSU_io_prf_0_idx[5:0]                                                     ), //o
    .io_prf_0_data                             (cpuClockingArea_prf_io_read_4_0_data[31:0]                                                                 ), //i
    .io_prf_1_idx                              (cpuClockingArea_areaFlushReset_roLSU_io_prf_1_idx[5:0]                                                     ), //o
    .io_prf_1_data                             (cpuClockingArea_prf_io_read_4_1_data[31:0]                                                                 ), //i
    .io_interrupt                              (cpuClockingArea_csr_io_interrupt                                                                           )  //i
  );
  ALU cpuClockingArea_areaFlushReset_fuALU0 (
    .io_input_valid                              (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_valid                             ), //i
    .io_input_ready                              (cpuClockingArea_areaFlushReset_fuALU0_io_input_ready                                             ), //o
    .io_input_payload_src1                       (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src1[31:0]                ), //i
    .io_input_payload_src2                       (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src2[31:0]                ), //i
    .io_input_payload_src3                       (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src3[31:0]                ), //i
    .io_input_payload_src4                       (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src4[31:0]                ), //i
    .io_input_payload_robIdx                     (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_robIdx[4:0]               ), //i
    .io_input_payload_branchInfo_predictPC       (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_branchInfo_predictPC[31:0]), //i
    .io_input_payload_branchInfo_predictResult   (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_branchInfo_predictResult  ), //i
    .io_input_payload_exceptionInfo_exception    (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_exceptionInfo_exception   ), //i
    .io_input_payload_exceptionInfo_eCode        (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_exceptionInfo_eCode[5:0]  ), //i
    .io_input_payload_exceptionInfo_eSubCode     (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode    ), //i
    .io_input_payload_pc                         (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_pc[31:0]                  ), //i
    .io_input_payload_prd                        (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_prd[5:0]                  ), //i
    .io_input_payload_uop_aluOp                  (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp[3:0]            ), //i
    .io_input_payload_uop_bruOp                  (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_bruOp[1:0]            ), //i
    .io_input_payload_uop_cruOp                  (toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_cruOp[1:0]            ), //i
    .io_output_valid                             (cpuClockingArea_areaFlushReset_fuALU0_io_output_valid                                            ), //o
    .io_output_ready                             (cpuClockingArea_areaFlushReset_fuALU0_io_output_ready                                            ), //i
    .io_output_payload_robIdx                    (cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_robIdx[4:0]                              ), //o
    .io_output_payload_data                      (cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_data[31:0]                               ), //o
    .io_output_payload_prd                       (cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_prd[5:0]                                 ), //o
    .io_output_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_branchResult_targetPC[31:0]              ), //o
    .io_output_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_branchResult_branchResult                ), //o
    .io_output_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_branchResult_predictFail                 ), //o
    .io_output_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_exceptionInfo_exception                  ), //o
    .io_output_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_exceptionInfo_eCode[5:0]                 ), //o
    .io_output_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_exceptionInfo_eSubCode                   ), //o
    .io_forward_valid                            (cpuClockingArea_areaFlushReset_fuALU0_io_forward_valid                                           ), //o
    .io_forward_payload_idx                      (cpuClockingArea_areaFlushReset_fuALU0_io_forward_payload_idx[5:0]                                ), //o
    .io_forward_payload_payload                  (cpuClockingArea_areaFlushReset_fuALU0_io_forward_payload_payload[31:0]                           ), //o
    .io_wakeOut_valid                            (cpuClockingArea_areaFlushReset_fuALU0_io_wakeOut_valid                                           ), //o
    .io_wakeOut_payload                          (cpuClockingArea_areaFlushReset_fuALU0_io_wakeOut_payload[5:0]                                    ), //o
    .io_csrWrite_value                           (cpuClockingArea_areaFlushReset_fuALU0_io_csrWrite_value[31:0]                                    ), //o
    .io_csrWrite_address                         (cpuClockingArea_areaFlushReset_fuALU0_io_csrWrite_address[13:0]                                  ), //o
    .io_csrWrite_wen                             (cpuClockingArea_areaFlushReset_fuALU0_io_csrWrite_wen                                            )  //o
  );
  ALU_1 cpuClockingArea_areaFlushReset_fuALU1 (
    .io_input_valid                              (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_valid                             ), //i
    .io_input_ready                              (cpuClockingArea_areaFlushReset_fuALU1_io_input_ready                                             ), //o
    .io_input_payload_src1                       (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src1[31:0]                ), //i
    .io_input_payload_src2                       (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src2[31:0]                ), //i
    .io_input_payload_src3                       (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src3[31:0]                ), //i
    .io_input_payload_src4                       (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src4[31:0]                ), //i
    .io_input_payload_robIdx                     (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_robIdx[4:0]               ), //i
    .io_input_payload_branchInfo_predictPC       (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_branchInfo_predictPC[31:0]), //i
    .io_input_payload_branchInfo_predictResult   (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_branchInfo_predictResult  ), //i
    .io_input_payload_exceptionInfo_exception    (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_exceptionInfo_exception   ), //i
    .io_input_payload_exceptionInfo_eCode        (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_exceptionInfo_eCode[5:0]  ), //i
    .io_input_payload_exceptionInfo_eSubCode     (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode    ), //i
    .io_input_payload_pc                         (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_pc[31:0]                  ), //i
    .io_input_payload_prd                        (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_prd[5:0]                  ), //i
    .io_input_payload_uop_aluOp                  (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp[3:0]            ), //i
    .io_input_payload_uop_bruOp                  (toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_bruOp[1:0]            ), //i
    .io_output_valid                             (cpuClockingArea_areaFlushReset_fuALU1_io_output_valid                                            ), //o
    .io_output_ready                             (cpuClockingArea_areaFlushReset_fuALU1_io_output_ready                                            ), //i
    .io_output_payload_robIdx                    (cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_robIdx[4:0]                              ), //o
    .io_output_payload_data                      (cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_data[31:0]                               ), //o
    .io_output_payload_prd                       (cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_prd[5:0]                                 ), //o
    .io_output_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_branchResult_targetPC[31:0]              ), //o
    .io_output_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_branchResult_branchResult                ), //o
    .io_output_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_branchResult_predictFail                 ), //o
    .io_output_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_exceptionInfo_exception                  ), //o
    .io_output_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_exceptionInfo_eCode[5:0]                 ), //o
    .io_output_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_exceptionInfo_eSubCode                   ), //o
    .io_forward_valid                            (cpuClockingArea_areaFlushReset_fuALU1_io_forward_valid                                           ), //o
    .io_forward_payload_idx                      (cpuClockingArea_areaFlushReset_fuALU1_io_forward_payload_idx[5:0]                                ), //o
    .io_forward_payload_payload                  (cpuClockingArea_areaFlushReset_fuALU1_io_forward_payload_payload[31:0]                           ), //o
    .io_wakeOut_valid                            (cpuClockingArea_areaFlushReset_fuALU1_io_wakeOut_valid                                           ), //o
    .io_wakeOut_payload                          (cpuClockingArea_areaFlushReset_fuALU1_io_wakeOut_payload[5:0]                                    )  //o
  );
  MULU cpuClockingArea_areaFlushReset_fuMULU (
    .io_input_valid                              (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_valid                              ), //i
    .io_input_ready                              (cpuClockingArea_areaFlushReset_fuMULU_io_input_ready                                              ), //o
    .io_input_payload_src1                       (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_src1[31:0]                 ), //i
    .io_input_payload_src2                       (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_src2[31:0]                 ), //i
    .io_input_payload_robIdx                     (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_robIdx[4:0]                ), //i
    .io_input_payload_branchResult_targetPC      (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_branchResult_targetPC[31:0]), //i
    .io_input_payload_branchResult_branchResult  (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_branchResult_branchResult  ), //i
    .io_input_payload_branchResult_predictFail   (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_branchResult_predictFail   ), //i
    .io_input_payload_exceptionInfo_exception    (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_exceptionInfo_exception    ), //i
    .io_input_payload_exceptionInfo_eCode        (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_exceptionInfo_eCode[5:0]   ), //i
    .io_input_payload_exceptionInfo_eSubCode     (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode     ), //i
    .io_input_payload_pc                         (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_pc[31:0]                   ), //i
    .io_input_payload_prd                        (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_prd[5:0]                   ), //i
    .io_input_payload_uop_muluOp                 (toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_uop_muluOp[1:0]            ), //i
    .io_output_valid                             (cpuClockingArea_areaFlushReset_fuMULU_io_output_valid                                             ), //o
    .io_output_ready                             (cpuClockingArea_areaFlushReset_fuMULU_io_output_ready                                             ), //i
    .io_output_payload_robIdx                    (cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_robIdx[4:0]                               ), //o
    .io_output_payload_data                      (cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_data[31:0]                                ), //o
    .io_output_payload_prd                       (cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_prd[5:0]                                  ), //o
    .io_output_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_branchResult_targetPC[31:0]               ), //o
    .io_output_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_branchResult_branchResult                 ), //o
    .io_output_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_branchResult_predictFail                  ), //o
    .io_output_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_exceptionInfo_exception                   ), //o
    .io_output_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_exceptionInfo_eCode[5:0]                  ), //o
    .io_output_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_exceptionInfo_eSubCode                    ), //o
    .io_forward_valid                            (cpuClockingArea_areaFlushReset_fuMULU_io_forward_valid                                            ), //o
    .io_forward_payload_idx                      (cpuClockingArea_areaFlushReset_fuMULU_io_forward_payload_idx[5:0]                                 ), //o
    .io_forward_payload_payload                  (cpuClockingArea_areaFlushReset_fuMULU_io_forward_payload_payload[31:0]                            ), //o
    .io_wakeOut_0_valid                          (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_0_valid                                          ), //o
    .io_wakeOut_0_payload                        (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_0_payload[5:0]                                   ), //o
    .io_wakeOut_1_valid                          (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_1_valid                                          ), //o
    .io_wakeOut_1_payload                        (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_1_payload[5:0]                                   ), //o
    .io_wakeOut_2_valid                          (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_2_valid                                          ), //o
    .io_wakeOut_2_payload                        (cpuClockingArea_areaFlushReset_fuMULU_io_wakeOut_2_payload[5:0]                                   ), //o
    .aclk                                        (aclk                                                                                              ), //i
    .cpuClockingArea_areaFlushReset_newReset     (cpuClockingArea_areaFlushReset_newReset                                                           )  //i
  );
  DIVU cpuClockingArea_areaFlushReset_fuDIVU (
    .io_input_valid                              (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_valid                              ), //i
    .io_input_ready                              (cpuClockingArea_areaFlushReset_fuDIVU_io_input_ready                                              ), //o
    .io_input_payload_src1                       (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_src1[31:0]                 ), //i
    .io_input_payload_src2                       (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_src2[31:0]                 ), //i
    .io_input_payload_robIdx                     (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_robIdx[4:0]                ), //i
    .io_input_payload_branchResult_targetPC      (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_branchResult_targetPC[31:0]), //i
    .io_input_payload_branchResult_branchResult  (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_branchResult_branchResult  ), //i
    .io_input_payload_branchResult_predictFail   (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_branchResult_predictFail   ), //i
    .io_input_payload_exceptionInfo_exception    (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_exceptionInfo_exception    ), //i
    .io_input_payload_exceptionInfo_eCode        (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_exceptionInfo_eCode[5:0]   ), //i
    .io_input_payload_exceptionInfo_eSubCode     (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode     ), //i
    .io_input_payload_pc                         (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_pc[31:0]                   ), //i
    .io_input_payload_prd                        (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_prd[5:0]                   ), //i
    .io_input_payload_uop_divuOp                 (toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_uop_divuOp[1:0]            ), //i
    .io_output_valid                             (cpuClockingArea_areaFlushReset_fuDIVU_io_output_valid                                             ), //o
    .io_output_ready                             (cpuClockingArea_areaFlushReset_fuDIVU_io_output_ready                                             ), //i
    .io_output_payload_robIdx                    (cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_robIdx[4:0]                               ), //o
    .io_output_payload_data                      (cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_data[31:0]                                ), //o
    .io_output_payload_prd                       (cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_prd[5:0]                                  ), //o
    .io_output_payload_branchResult_targetPC     (cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_branchResult_targetPC[31:0]               ), //o
    .io_output_payload_branchResult_branchResult (cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_branchResult_branchResult                 ), //o
    .io_output_payload_branchResult_predictFail  (cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_branchResult_predictFail                  ), //o
    .io_output_payload_exceptionInfo_exception   (cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_exceptionInfo_exception                   ), //o
    .io_output_payload_exceptionInfo_eCode       (cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_exceptionInfo_eCode[5:0]                  ), //o
    .io_output_payload_exceptionInfo_eSubCode    (cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_exceptionInfo_eSubCode                    ), //o
    .aclk                                        (aclk                                                                                              ), //i
    .cpuClockingArea_areaFlushReset_newReset     (cpuClockingArea_areaFlushReset_newReset                                                           )  //i
  );
  CommitLogic cpuClockingArea_areaFlushReset_commitALU0 (
    .io_input_valid                             (toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_valid                              ), //i
    .io_input_ready                             (cpuClockingArea_areaFlushReset_commitALU0_io_input_ready                                            ), //o
    .io_input_payload_robIdx                    (toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_robIdx[4:0]                ), //i
    .io_input_payload_data                      (toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_data[31:0]                 ), //i
    .io_input_payload_prd                       (toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_prd[5:0]                   ), //i
    .io_input_payload_branchResult_targetPC     (toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_branchResult_targetPC[31:0]), //i
    .io_input_payload_branchResult_branchResult (toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_branchResult_branchResult  ), //i
    .io_input_payload_branchResult_predictFail  (toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_branchResult_predictFail   ), //i
    .io_input_payload_exceptionInfo_exception   (toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_exceptionInfo_exception    ), //i
    .io_input_payload_exceptionInfo_eCode       (toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_exceptionInfo_eCode[5:0]   ), //i
    .io_input_payload_exceptionInfo_eSubCode    (toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_exceptionInfo_eSubCode     ), //i
    .io_srat_prd                                (cpuClockingArea_areaFlushReset_commitALU0_io_srat_prd[5:0]                                          ), //o
    .io_srat_wen                                (cpuClockingArea_areaFlushReset_commitALU0_io_srat_wen                                               ), //o
    .io_rob_robIdx                              (cpuClockingArea_areaFlushReset_commitALU0_io_rob_robIdx[4:0]                                        ), //o
    .io_rob_branchResult_targetPC               (cpuClockingArea_areaFlushReset_commitALU0_io_rob_branchResult_targetPC[31:0]                        ), //o
    .io_rob_branchResult_branchResult           (cpuClockingArea_areaFlushReset_commitALU0_io_rob_branchResult_branchResult                          ), //o
    .io_rob_branchResult_predictFail            (cpuClockingArea_areaFlushReset_commitALU0_io_rob_branchResult_predictFail                           ), //o
    .io_rob_exceptionInfo_exception             (cpuClockingArea_areaFlushReset_commitALU0_io_rob_exceptionInfo_exception                            ), //o
    .io_rob_exceptionInfo_eCode                 (cpuClockingArea_areaFlushReset_commitALU0_io_rob_exceptionInfo_eCode[5:0]                           ), //o
    .io_rob_exceptionInfo_eSubCode              (cpuClockingArea_areaFlushReset_commitALU0_io_rob_exceptionInfo_eSubCode                             ), //o
    .io_rob_valid                               (cpuClockingArea_areaFlushReset_commitALU0_io_rob_valid                                              ), //o
    .io_prf_idx                                 (cpuClockingArea_areaFlushReset_commitALU0_io_prf_idx[5:0]                                           ), //o
    .io_prf_data                                (cpuClockingArea_areaFlushReset_commitALU0_io_prf_data[31:0]                                         ), //o
    .io_forward_valid                           (cpuClockingArea_areaFlushReset_commitALU0_io_forward_valid                                          ), //o
    .io_forward_payload_idx                     (cpuClockingArea_areaFlushReset_commitALU0_io_forward_payload_idx[5:0]                               ), //o
    .io_forward_payload_payload                 (cpuClockingArea_areaFlushReset_commitALU0_io_forward_payload_payload[31:0]                          )  //o
  );
  CommitLogic cpuClockingArea_areaFlushReset_commitALU1 (
    .io_input_valid                             (toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_valid                              ), //i
    .io_input_ready                             (cpuClockingArea_areaFlushReset_commitALU1_io_input_ready                                            ), //o
    .io_input_payload_robIdx                    (toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_robIdx[4:0]                ), //i
    .io_input_payload_data                      (toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_data[31:0]                 ), //i
    .io_input_payload_prd                       (toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_prd[5:0]                   ), //i
    .io_input_payload_branchResult_targetPC     (toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_branchResult_targetPC[31:0]), //i
    .io_input_payload_branchResult_branchResult (toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_branchResult_branchResult  ), //i
    .io_input_payload_branchResult_predictFail  (toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_branchResult_predictFail   ), //i
    .io_input_payload_exceptionInfo_exception   (toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_exceptionInfo_exception    ), //i
    .io_input_payload_exceptionInfo_eCode       (toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_exceptionInfo_eCode[5:0]   ), //i
    .io_input_payload_exceptionInfo_eSubCode    (toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_exceptionInfo_eSubCode     ), //i
    .io_srat_prd                                (cpuClockingArea_areaFlushReset_commitALU1_io_srat_prd[5:0]                                          ), //o
    .io_srat_wen                                (cpuClockingArea_areaFlushReset_commitALU1_io_srat_wen                                               ), //o
    .io_rob_robIdx                              (cpuClockingArea_areaFlushReset_commitALU1_io_rob_robIdx[4:0]                                        ), //o
    .io_rob_branchResult_targetPC               (cpuClockingArea_areaFlushReset_commitALU1_io_rob_branchResult_targetPC[31:0]                        ), //o
    .io_rob_branchResult_branchResult           (cpuClockingArea_areaFlushReset_commitALU1_io_rob_branchResult_branchResult                          ), //o
    .io_rob_branchResult_predictFail            (cpuClockingArea_areaFlushReset_commitALU1_io_rob_branchResult_predictFail                           ), //o
    .io_rob_exceptionInfo_exception             (cpuClockingArea_areaFlushReset_commitALU1_io_rob_exceptionInfo_exception                            ), //o
    .io_rob_exceptionInfo_eCode                 (cpuClockingArea_areaFlushReset_commitALU1_io_rob_exceptionInfo_eCode[5:0]                           ), //o
    .io_rob_exceptionInfo_eSubCode              (cpuClockingArea_areaFlushReset_commitALU1_io_rob_exceptionInfo_eSubCode                             ), //o
    .io_rob_valid                               (cpuClockingArea_areaFlushReset_commitALU1_io_rob_valid                                              ), //o
    .io_prf_idx                                 (cpuClockingArea_areaFlushReset_commitALU1_io_prf_idx[5:0]                                           ), //o
    .io_prf_data                                (cpuClockingArea_areaFlushReset_commitALU1_io_prf_data[31:0]                                         ), //o
    .io_forward_valid                           (cpuClockingArea_areaFlushReset_commitALU1_io_forward_valid                                          ), //o
    .io_forward_payload_idx                     (cpuClockingArea_areaFlushReset_commitALU1_io_forward_payload_idx[5:0]                               ), //o
    .io_forward_payload_payload                 (cpuClockingArea_areaFlushReset_commitALU1_io_forward_payload_payload[31:0]                          )  //o
  );
  CommitLogic cpuClockingArea_areaFlushReset_commitMULU (
    .io_input_valid                             (toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_valid                              ), //i
    .io_input_ready                             (cpuClockingArea_areaFlushReset_commitMULU_io_input_ready                                            ), //o
    .io_input_payload_robIdx                    (toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_robIdx[4:0]                ), //i
    .io_input_payload_data                      (toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_data[31:0]                 ), //i
    .io_input_payload_prd                       (toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_prd[5:0]                   ), //i
    .io_input_payload_branchResult_targetPC     (toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_branchResult_targetPC[31:0]), //i
    .io_input_payload_branchResult_branchResult (toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_branchResult_branchResult  ), //i
    .io_input_payload_branchResult_predictFail  (toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_branchResult_predictFail   ), //i
    .io_input_payload_exceptionInfo_exception   (toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_exceptionInfo_exception    ), //i
    .io_input_payload_exceptionInfo_eCode       (toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_exceptionInfo_eCode[5:0]   ), //i
    .io_input_payload_exceptionInfo_eSubCode    (toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_exceptionInfo_eSubCode     ), //i
    .io_srat_prd                                (cpuClockingArea_areaFlushReset_commitMULU_io_srat_prd[5:0]                                          ), //o
    .io_srat_wen                                (cpuClockingArea_areaFlushReset_commitMULU_io_srat_wen                                               ), //o
    .io_rob_robIdx                              (cpuClockingArea_areaFlushReset_commitMULU_io_rob_robIdx[4:0]                                        ), //o
    .io_rob_branchResult_targetPC               (cpuClockingArea_areaFlushReset_commitMULU_io_rob_branchResult_targetPC[31:0]                        ), //o
    .io_rob_branchResult_branchResult           (cpuClockingArea_areaFlushReset_commitMULU_io_rob_branchResult_branchResult                          ), //o
    .io_rob_branchResult_predictFail            (cpuClockingArea_areaFlushReset_commitMULU_io_rob_branchResult_predictFail                           ), //o
    .io_rob_exceptionInfo_exception             (cpuClockingArea_areaFlushReset_commitMULU_io_rob_exceptionInfo_exception                            ), //o
    .io_rob_exceptionInfo_eCode                 (cpuClockingArea_areaFlushReset_commitMULU_io_rob_exceptionInfo_eCode[5:0]                           ), //o
    .io_rob_exceptionInfo_eSubCode              (cpuClockingArea_areaFlushReset_commitMULU_io_rob_exceptionInfo_eSubCode                             ), //o
    .io_rob_valid                               (cpuClockingArea_areaFlushReset_commitMULU_io_rob_valid                                              ), //o
    .io_prf_idx                                 (cpuClockingArea_areaFlushReset_commitMULU_io_prf_idx[5:0]                                           ), //o
    .io_prf_data                                (cpuClockingArea_areaFlushReset_commitMULU_io_prf_data[31:0]                                         ), //o
    .io_forward_valid                           (cpuClockingArea_areaFlushReset_commitMULU_io_forward_valid                                          ), //o
    .io_forward_payload_idx                     (cpuClockingArea_areaFlushReset_commitMULU_io_forward_payload_idx[5:0]                               ), //o
    .io_forward_payload_payload                 (cpuClockingArea_areaFlushReset_commitMULU_io_forward_payload_payload[31:0]                          )  //o
  );
  CommitLogic cpuClockingArea_areaFlushReset_commitDIVU (
    .io_input_valid                             (toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_valid                              ), //i
    .io_input_ready                             (cpuClockingArea_areaFlushReset_commitDIVU_io_input_ready                                            ), //o
    .io_input_payload_robIdx                    (toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_robIdx[4:0]                ), //i
    .io_input_payload_data                      (toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_data[31:0]                 ), //i
    .io_input_payload_prd                       (toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_prd[5:0]                   ), //i
    .io_input_payload_branchResult_targetPC     (toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_branchResult_targetPC[31:0]), //i
    .io_input_payload_branchResult_branchResult (toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_branchResult_branchResult  ), //i
    .io_input_payload_branchResult_predictFail  (toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_branchResult_predictFail   ), //i
    .io_input_payload_exceptionInfo_exception   (toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_exceptionInfo_exception    ), //i
    .io_input_payload_exceptionInfo_eCode       (toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_exceptionInfo_eCode[5:0]   ), //i
    .io_input_payload_exceptionInfo_eSubCode    (toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_exceptionInfo_eSubCode     ), //i
    .io_srat_prd                                (cpuClockingArea_areaFlushReset_commitDIVU_io_srat_prd[5:0]                                          ), //o
    .io_srat_wen                                (cpuClockingArea_areaFlushReset_commitDIVU_io_srat_wen                                               ), //o
    .io_rob_robIdx                              (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_robIdx[4:0]                                        ), //o
    .io_rob_branchResult_targetPC               (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_branchResult_targetPC[31:0]                        ), //o
    .io_rob_branchResult_branchResult           (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_branchResult_branchResult                          ), //o
    .io_rob_branchResult_predictFail            (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_branchResult_predictFail                           ), //o
    .io_rob_exceptionInfo_exception             (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_exceptionInfo_exception                            ), //o
    .io_rob_exceptionInfo_eCode                 (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_exceptionInfo_eCode[5:0]                           ), //o
    .io_rob_exceptionInfo_eSubCode              (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_exceptionInfo_eSubCode                             ), //o
    .io_rob_valid                               (cpuClockingArea_areaFlushReset_commitDIVU_io_rob_valid                                              ), //o
    .io_prf_idx                                 (cpuClockingArea_areaFlushReset_commitDIVU_io_prf_idx[5:0]                                           ), //o
    .io_prf_data                                (cpuClockingArea_areaFlushReset_commitDIVU_io_prf_data[31:0]                                         ), //o
    .io_forward_valid                           (cpuClockingArea_areaFlushReset_commitDIVU_io_forward_valid                                          ), //o
    .io_forward_payload_idx                     (cpuClockingArea_areaFlushReset_commitDIVU_io_forward_payload_idx[5:0]                               ), //o
    .io_forward_payload_payload                 (cpuClockingArea_areaFlushReset_commitDIVU_io_forward_payload_payload[31:0]                          )  //o
  );
  CommitLogic cpuClockingArea_areaFlushReset_commitLSU (
    .io_input_valid                             (toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_valid                              ), //i
    .io_input_ready                             (cpuClockingArea_areaFlushReset_commitLSU_io_input_ready                             ), //o
    .io_input_payload_robIdx                    (toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_robIdx[4:0]                ), //i
    .io_input_payload_data                      (toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_data[31:0]                 ), //i
    .io_input_payload_prd                       (toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_prd[5:0]                   ), //i
    .io_input_payload_branchResult_targetPC     (toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_branchResult_targetPC[31:0]), //i
    .io_input_payload_branchResult_branchResult (toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_branchResult_branchResult  ), //i
    .io_input_payload_branchResult_predictFail  (toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_branchResult_predictFail   ), //i
    .io_input_payload_exceptionInfo_exception   (toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_exceptionInfo_exception    ), //i
    .io_input_payload_exceptionInfo_eCode       (toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_exceptionInfo_eCode[5:0]   ), //i
    .io_input_payload_exceptionInfo_eSubCode    (toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_exceptionInfo_eSubCode     ), //i
    .io_srat_prd                                (cpuClockingArea_areaFlushReset_commitLSU_io_srat_prd[5:0]                           ), //o
    .io_srat_wen                                (cpuClockingArea_areaFlushReset_commitLSU_io_srat_wen                                ), //o
    .io_rob_robIdx                              (cpuClockingArea_areaFlushReset_commitLSU_io_rob_robIdx[4:0]                         ), //o
    .io_rob_branchResult_targetPC               (cpuClockingArea_areaFlushReset_commitLSU_io_rob_branchResult_targetPC[31:0]         ), //o
    .io_rob_branchResult_branchResult           (cpuClockingArea_areaFlushReset_commitLSU_io_rob_branchResult_branchResult           ), //o
    .io_rob_branchResult_predictFail            (cpuClockingArea_areaFlushReset_commitLSU_io_rob_branchResult_predictFail            ), //o
    .io_rob_exceptionInfo_exception             (cpuClockingArea_areaFlushReset_commitLSU_io_rob_exceptionInfo_exception             ), //o
    .io_rob_exceptionInfo_eCode                 (cpuClockingArea_areaFlushReset_commitLSU_io_rob_exceptionInfo_eCode[5:0]            ), //o
    .io_rob_exceptionInfo_eSubCode              (cpuClockingArea_areaFlushReset_commitLSU_io_rob_exceptionInfo_eSubCode              ), //o
    .io_rob_valid                               (cpuClockingArea_areaFlushReset_commitLSU_io_rob_valid                               ), //o
    .io_prf_idx                                 (cpuClockingArea_areaFlushReset_commitLSU_io_prf_idx[5:0]                            ), //o
    .io_prf_data                                (cpuClockingArea_areaFlushReset_commitLSU_io_prf_data[31:0]                          ), //o
    .io_forward_valid                           (cpuClockingArea_areaFlushReset_commitLSU_io_forward_valid                           ), //o
    .io_forward_payload_idx                     (cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_idx[5:0]                ), //o
    .io_forward_payload_payload                 (cpuClockingArea_areaFlushReset_commitLSU_io_forward_payload_payload[31:0]           )  //o
  );
  always @(*) begin
    case(_zz_DaRAT_val_1_1)
      6'b000000 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_1 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_2_1)
      6'b000000 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_2 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_3_1)
      6'b000000 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_3 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_4_1)
      6'b000000 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_4 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_5_1)
      6'b000000 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_5 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_6_1)
      6'b000000 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_6 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_7_1)
      6'b000000 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_7 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_8_1)
      6'b000000 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_8 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_9_1)
      6'b000000 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_9 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_10_1)
      6'b000000 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_10 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_11_1)
      6'b000000 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_11 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_12_1)
      6'b000000 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_12 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_13_1)
      6'b000000 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_13 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_14_1)
      6'b000000 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_14 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_15_1)
      6'b000000 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_15 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_16_1)
      6'b000000 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_16 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_17_1)
      6'b000000 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_17 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_18_1)
      6'b000000 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_18 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_19_1)
      6'b000000 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_19 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_20_1)
      6'b000000 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_20 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_21_1)
      6'b000000 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_21 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_22_1)
      6'b000000 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_22 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_23_1)
      6'b000000 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_23 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_24_1)
      6'b000000 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_24 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_25_1)
      6'b000000 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_25 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_26_1)
      6'b000000 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_26 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_27_1)
      6'b000000 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_27 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_28_1)
      6'b000000 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_28 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_29_1)
      6'b000000 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_29 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_30_1)
      6'b000000 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_30 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  always @(*) begin
    case(_zz_DaRAT_val_31_1)
      6'b000000 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_0;
      6'b000001 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_1;
      6'b000010 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_2;
      6'b000011 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_3;
      6'b000100 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_4;
      6'b000101 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_5;
      6'b000110 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_6;
      6'b000111 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_7;
      6'b001000 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_8;
      6'b001001 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_9;
      6'b001010 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_10;
      6'b001011 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_11;
      6'b001100 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_12;
      6'b001101 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_13;
      6'b001110 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_14;
      6'b001111 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_15;
      6'b010000 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_16;
      6'b010001 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_17;
      6'b010010 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_18;
      6'b010011 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_19;
      6'b010100 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_20;
      6'b010101 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_21;
      6'b010110 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_22;
      6'b010111 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_23;
      6'b011000 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_24;
      6'b011001 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_25;
      6'b011010 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_26;
      6'b011011 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_27;
      6'b011100 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_28;
      6'b011101 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_29;
      6'b011110 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_30;
      6'b011111 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_31;
      6'b100000 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_32;
      6'b100001 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_33;
      6'b100010 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_34;
      6'b100011 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_35;
      6'b100100 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_36;
      6'b100101 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_37;
      6'b100110 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_38;
      6'b100111 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_39;
      6'b101000 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_40;
      6'b101001 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_41;
      6'b101010 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_42;
      6'b101011 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_43;
      6'b101100 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_44;
      6'b101101 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_45;
      6'b101110 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_46;
      6'b101111 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_47;
      6'b110000 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_48;
      6'b110001 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_49;
      6'b110010 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_50;
      6'b110011 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_51;
      6'b110100 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_52;
      6'b110101 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_53;
      6'b110110 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_54;
      6'b110111 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_55;
      6'b111000 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_56;
      6'b111001 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_57;
      6'b111010 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_58;
      6'b111011 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_59;
      6'b111100 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_60;
      6'b111101 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_61;
      6'b111110 : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_62;
      default : _zz_DaRAT_val_31 = cpuClockingArea_prf_io_debugRegs_63;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp)
      ALUOp_add : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "passa";
      ALUOp_passb : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "passb";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_bruOp)
      BRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_bruOp_string = "ncadd";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_cruOp)
      CRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_cruOp_string = "nop ";
      CRUOp_pass : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_cruOp_string = "pass";
      CRUOp_mask : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_cruOp_string = "mask";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp)
      ALUROOp_reg_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp_string = "linkreg";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp)
      ALUOp_add : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "add  ";
      ALUOp_sub : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "sub  ";
      ALUOp_slt : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "slt  ";
      ALUOp_sltu : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "sltu ";
      ALUOp_eq : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "and_1";
      ALUOp_or_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "sra_1";
      ALUOp_passa : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "passa";
      ALUOp_passb : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "passb";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_bruOp)
      BRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_bruOp_string = "nop  ";
      BRUOp_add : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_bruOp_string = "add  ";
      BRUOp_cadd : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_bruOp_string = "ncadd";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_cruOp)
      CRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_cruOp_string = "nop ";
      CRUOp_pass : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_cruOp_string = "pass";
      CRUOp_mask : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_cruOp_string = "mask";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp)
      ALUROOp_reg_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp_string = "linkreg";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp)
      ALUOp_add : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "passa";
      ALUOp_passb : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "passb";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_bruOp)
      BRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_bruOp_string = "ncadd";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp)
      ALUROOp_reg_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp_string = "linkreg";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_cruROOp)
      CRUROOp_id : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_cruROOp_string = "id";
      CRUROOp_lo : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_cruROOp_string = "lo";
      CRUROOp_hi : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_cruROOp_string = "hi";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp)
      ALUOp_add : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "add  ";
      ALUOp_sub : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "sub  ";
      ALUOp_slt : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "slt  ";
      ALUOp_sltu : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "sltu ";
      ALUOp_eq : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "and_1";
      ALUOp_or_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "sra_1";
      ALUOp_passa : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "passa";
      ALUOp_passb : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "passb";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_bruOp)
      BRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_bruOp_string = "nop  ";
      BRUOp_add : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_bruOp_string = "add  ";
      BRUOp_cadd : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_bruOp_string = "ncadd";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp)
      ALUROOp_reg_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp_string = "linkreg";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_cruROOp)
      CRUROOp_id : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_cruROOp_string = "id";
      CRUROOp_lo : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_cruROOp_string = "lo";
      CRUROOp_hi : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_cruROOp_string = "hi";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_uop_muluOp)
      MULUOp_mullo : toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_uop_muluOp_string = "mulhiu";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_uop_muluOp)
      MULUOp_mullo : toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_uop_muluOp_string = "mulhiu";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_uop_divuOp)
      DIVUOp_div : toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_uop_divuOp_string = "div  ";
      DIVUOp_divu : toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_uop_divuOp_string = "mod_1";
      DIVUOp_modu : toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_uop_divuOp_string = "modu ";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_uop_divuOp)
      DIVUOp_div : toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_uop_divuOp_string = "div  ";
      DIVUOp_divu : toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_uop_divuOp_string = "mod_1";
      DIVUOp_modu : toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_uop_divuOp_string = "modu ";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp)
      LSUOp_cacop : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "ll     ";
      LSUOp_sc : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "sc     ";
      LSUOp_ld : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "ldu    ";
      LSUOp_st : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "st     ";
      LSUOp_preld : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "ibar   ";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_roop_lsuROOp)
      LSUROOp_reg_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_roop_lsuROOp_string = "regimm";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp)
      LSUOp_cacop : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "ll     ";
      LSUOp_sc : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "sc     ";
      LSUOp_ld : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "ldu    ";
      LSUOp_st : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "st     ";
      LSUOp_preld : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "ibar   ";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_roop_lsuROOp)
      LSUROOp_reg_1 : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_roop_lsuROOp_string = "regimm";
      default : toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp)
      ALUOp_add : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "passa";
      ALUOp_passb : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "passb";
      default : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_bruOp)
      BRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_bruOp_string = "ncadd";
      default : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_cruOp)
      CRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_cruOp_string = "nop ";
      CRUOp_pass : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_cruOp_string = "pass";
      CRUOp_mask : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_cruOp_string = "mask";
      default : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp)
      ALUOp_add : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "add  ";
      ALUOp_sub : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "sub  ";
      ALUOp_slt : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "slt  ";
      ALUOp_sltu : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "sltu ";
      ALUOp_eq : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "and_1";
      ALUOp_or_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "sra_1";
      ALUOp_passa : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "passa";
      ALUOp_passb : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "passb";
      default : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_bruOp)
      BRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_bruOp_string = "nop  ";
      BRUOp_add : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_bruOp_string = "add  ";
      BRUOp_cadd : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_bruOp_string = "ncadd";
      default : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_cruOp)
      CRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_cruOp_string = "nop ";
      CRUOp_pass : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_cruOp_string = "pass";
      CRUOp_mask : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_cruOp_string = "mask";
      default : toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp)
      ALUOp_add : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "passa";
      ALUOp_passb : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "passb";
      default : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_bruOp)
      BRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_bruOp_string = "ncadd";
      default : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp)
      ALUOp_add : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "add  ";
      ALUOp_sub : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "sub  ";
      ALUOp_slt : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "slt  ";
      ALUOp_sltu : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "sltu ";
      ALUOp_eq : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "and_1";
      ALUOp_or_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "sra_1";
      ALUOp_passa : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "passa";
      ALUOp_passb : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "passb";
      default : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_bruOp)
      BRUOp_nop : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_bruOp_string = "nop  ";
      BRUOp_add : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_bruOp_string = "add  ";
      BRUOp_cadd : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_bruOp_string = "ncadd";
      default : toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_uop_muluOp)
      MULUOp_mullo : toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_uop_muluOp_string = "mulhiu";
      default : toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_uop_muluOp)
      MULUOp_mullo : toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_uop_muluOp_string = "mulhiu";
      default : toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_uop_divuOp)
      DIVUOp_div : toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_uop_divuOp_string = "div  ";
      DIVUOp_divu : toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_uop_divuOp_string = "mod_1";
      DIVUOp_modu : toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_uop_divuOp_string = "modu ";
      default : toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_uop_divuOp)
      DIVUOp_div : toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_uop_divuOp_string = "div  ";
      DIVUOp_divu : toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_uop_divuOp_string = "mod_1";
      DIVUOp_modu : toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_uop_divuOp_string = "modu ";
      default : toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp)
      LSUOp_cacop : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "ll     ";
      LSUOp_sc : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "sc     ";
      LSUOp_ld : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "ldu    ";
      LSUOp_st : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "st     ";
      LSUOp_preld : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "ibar   ";
      default : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp)
      LSUOp_cacop : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "ll     ";
      LSUOp_sc : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "sc     ";
      LSUOp_ld : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "ldu    ";
      LSUOp_st : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "st     ";
      LSUOp_preld : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "ibar   ";
      default : toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp_string = "???????";
    endcase
  end
  `endif

  assign DifftestBundle_DifftestTrapEventValid = 1'b0;
  assign cpuClockingArea_areaFlushReset_newReset = (aresetn && (! cpuClockingArea_rob_io_flush));
  always @(*) begin
    cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_ready = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_ready;
    if(when_Stream_l369) begin
      cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l369 = (! toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_branchInfo_predictPC = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_branchInfo_predictPC;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_branchInfo_predictResult = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_branchInfo_predictResult;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_pc = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_pc;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_psrc_0 = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_psrc_0;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_psrc_1 = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_psrc_1;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_imm = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_imm;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_aluOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_bruOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_bruOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_uop_cruOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_cruOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_payload_roop_aluROOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_m2sPipe_ready = cpuClockingArea_areaFlushReset_roALU0_io_cmd_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_ready = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_ready;
    if(when_Stream_l369_1) begin
      cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l369_1 = (! toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_branchInfo_predictPC = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_branchInfo_predictPC;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_branchInfo_predictResult = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_branchInfo_predictResult;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_pc = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_pc;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_psrc_0 = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_psrc_0;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_psrc_1 = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_psrc_1;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_imm = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_imm;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_aluOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_uop_bruOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_bruOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_aluROOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_payload_roop_cruROOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_cruROOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_m2sPipe_ready = cpuClockingArea_areaFlushReset_roALU1_io_cmd_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_ready = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_ready;
    if(when_Stream_l369_2) begin
      cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l369_2 = (! toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_branchResult_targetPC = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_branchResult_targetPC;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_branchResult_branchResult = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_branchResult_branchResult;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_branchResult_predictFail = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_branchResult_predictFail;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_pc = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_pc;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_psrc_0 = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_psrc_0;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_psrc_1 = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_psrc_1;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_imm = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_imm;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_payload_uop_muluOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_uop_muluOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_m2sPipe_ready = cpuClockingArea_areaFlushReset_roMULU_io_cmd_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_ready = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_ready;
    if(when_Stream_l369_3) begin
      cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l369_3 = (! toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_branchResult_targetPC = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_branchResult_targetPC;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_branchResult_branchResult = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_branchResult_branchResult;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_branchResult_predictFail = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_branchResult_predictFail;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_pc = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_pc;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_psrc_0 = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_psrc_0;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_psrc_1 = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_psrc_1;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_imm = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_imm;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_payload_uop_divuOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_uop_divuOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_m2sPipe_ready = cpuClockingArea_areaFlushReset_roDIVU_io_cmd_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_ready = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_ready;
    if(when_Stream_l369_4) begin
      cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l369_4 = (! toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_branchResult_targetPC = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_branchResult_targetPC;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_branchResult_branchResult = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_branchResult_branchResult;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_branchResult_predictFail = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_branchResult_predictFail;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_pc = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_pc;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_psrc_0 = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_psrc_0;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_psrc_1 = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_psrc_1;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_imm = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_imm;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_uop_lsuCoOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuCoOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_payload_roop_lsuROOp = toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_roop_lsuROOp;
  assign toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_m2sPipe_ready = cpuClockingArea_areaFlushReset_roLSU_io_cmd_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_roALU0_io_toFU_ready = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_ready;
    if(when_Stream_l369_5) begin
      cpuClockingArea_areaFlushReset_roALU0_io_toFU_ready = 1'b1;
    end
  end

  assign when_Stream_l369_5 = (! toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src1 = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src1;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src2 = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src2;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src3 = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src3;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_src4 = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src4;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_branchInfo_predictPC = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_branchInfo_predictPC;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_branchInfo_predictResult = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_branchInfo_predictResult;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_pc = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_pc;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_aluOp = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_bruOp = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_bruOp;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_payload_uop_cruOp = toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_cruOp;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_m2sPipe_ready = cpuClockingArea_areaFlushReset_fuALU0_io_input_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_roALU1_io_toFU_ready = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_ready;
    if(when_Stream_l369_6) begin
      cpuClockingArea_areaFlushReset_roALU1_io_toFU_ready = 1'b1;
    end
  end

  assign when_Stream_l369_6 = (! toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src1 = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src1;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src2 = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src2;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src3 = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src3;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_src4 = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src4;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_branchInfo_predictPC = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_branchInfo_predictPC;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_branchInfo_predictResult = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_branchInfo_predictResult;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_pc = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_pc;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_aluOp = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_payload_uop_bruOp = toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_bruOp;
  assign toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_m2sPipe_ready = cpuClockingArea_areaFlushReset_fuALU1_io_input_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_roMULU_io_toFU_ready = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_ready;
    if(when_Stream_l369_7) begin
      cpuClockingArea_areaFlushReset_roMULU_io_toFU_ready = 1'b1;
    end
  end

  assign when_Stream_l369_7 = (! toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_src1 = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_src1;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_src2 = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_src2;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_branchResult_targetPC = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_branchResult_targetPC;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_branchResult_branchResult = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_branchResult_branchResult;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_branchResult_predictFail = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_branchResult_predictFail;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_pc = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_pc;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_payload_uop_muluOp = toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_uop_muluOp;
  assign toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_m2sPipe_ready = cpuClockingArea_areaFlushReset_fuMULU_io_input_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_roDIVU_io_toFU_ready = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_ready;
    if(when_Stream_l369_8) begin
      cpuClockingArea_areaFlushReset_roDIVU_io_toFU_ready = 1'b1;
    end
  end

  assign when_Stream_l369_8 = (! toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_src1 = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_src1;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_src2 = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_src2;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_branchResult_targetPC = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_branchResult_targetPC;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_branchResult_branchResult = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_branchResult_branchResult;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_branchResult_predictFail = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_branchResult_predictFail;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_pc = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_pc;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_payload_uop_divuOp = toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_uop_divuOp;
  assign toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_m2sPipe_ready = cpuClockingArea_areaFlushReset_fuDIVU_io_input_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_roLSU_io_toFU_ready = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_ready;
    if(when_Stream_l369_9) begin
      cpuClockingArea_areaFlushReset_roLSU_io_toFU_ready = 1'b1;
    end
  end

  assign when_Stream_l369_9 = (! toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_src1 = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_src1;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_src2 = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_src2;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_src3 = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_src3;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_branchResult_targetPC = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_branchResult_targetPC;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_branchResult_branchResult = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_branchResult_branchResult;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_branchResult_predictFail = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_branchResult_predictFail;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_pc = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_pc;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuOp = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_payload_uop_lsuCoOp = toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuCoOp;
  assign toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_m2sPipe_ready = cpuClockingArea_fuLSU_io_input_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_fuALU0_io_output_ready = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_ready;
    if(when_Stream_l369_10) begin
      cpuClockingArea_areaFlushReset_fuALU0_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l369_10 = (! toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_data = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_data;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_branchResult_targetPC = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_branchResult_targetPC;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_branchResult_branchResult = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_branchResult_branchResult;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_branchResult_predictFail = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_branchResult_predictFail;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_ready = cpuClockingArea_areaFlushReset_commitALU0_io_input_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_fuALU1_io_output_ready = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_ready;
    if(when_Stream_l369_11) begin
      cpuClockingArea_areaFlushReset_fuALU1_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l369_11 = (! toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_data = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_data;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_branchResult_targetPC = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_branchResult_targetPC;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_branchResult_branchResult = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_branchResult_branchResult;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_branchResult_predictFail = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_branchResult_predictFail;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_ready = cpuClockingArea_areaFlushReset_commitALU1_io_input_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_fuMULU_io_output_ready = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_ready;
    if(when_Stream_l369_12) begin
      cpuClockingArea_areaFlushReset_fuMULU_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l369_12 = (! toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_data = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_data;
  assign toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_branchResult_targetPC = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_branchResult_targetPC;
  assign toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_branchResult_branchResult = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_branchResult_branchResult;
  assign toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_branchResult_predictFail = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_branchResult_predictFail;
  assign toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_ready = cpuClockingArea_areaFlushReset_commitMULU_io_input_ready;
  always @(*) begin
    cpuClockingArea_areaFlushReset_fuDIVU_io_output_ready = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_ready;
    if(when_Stream_l369_13) begin
      cpuClockingArea_areaFlushReset_fuDIVU_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l369_13 = (! toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_valid);
  assign toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_valid = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rValid;
  assign toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_robIdx;
  assign toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_data = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_data;
  assign toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_prd = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_prd;
  assign toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_branchResult_targetPC = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_branchResult_targetPC;
  assign toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_branchResult_branchResult = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_branchResult_branchResult;
  assign toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_branchResult_predictFail = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_branchResult_predictFail;
  assign toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_ready = cpuClockingArea_areaFlushReset_commitDIVU_io_input_ready;
  always @(*) begin
    cpuClockingArea_fuLSU_io_output_ready = toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_ready;
    if(when_Stream_l369_14) begin
      cpuClockingArea_fuLSU_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l369_14 = (! toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_valid);
  assign toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_valid = toplevel_cpuClockingArea_fuLSU_io_output_rValid;
  assign toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_robIdx = toplevel_cpuClockingArea_fuLSU_io_output_rData_robIdx;
  assign toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_data = toplevel_cpuClockingArea_fuLSU_io_output_rData_data;
  assign toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_prd = toplevel_cpuClockingArea_fuLSU_io_output_rData_prd;
  assign toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_branchResult_targetPC = toplevel_cpuClockingArea_fuLSU_io_output_rData_branchResult_targetPC;
  assign toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_branchResult_branchResult = toplevel_cpuClockingArea_fuLSU_io_output_rData_branchResult_branchResult;
  assign toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_branchResult_predictFail = toplevel_cpuClockingArea_fuLSU_io_output_rData_branchResult_predictFail;
  assign toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_exceptionInfo_exception = toplevel_cpuClockingArea_fuLSU_io_output_rData_exceptionInfo_exception;
  assign toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_exceptionInfo_eCode = toplevel_cpuClockingArea_fuLSU_io_output_rData_exceptionInfo_eCode;
  assign toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_exceptionInfo_eSubCode = toplevel_cpuClockingArea_fuLSU_io_output_rData_exceptionInfo_eSubCode;
  assign toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_ready = cpuClockingArea_areaFlushReset_commitLSU_io_input_ready;
  assign DaRAT_val_1 = _zz_DaRAT_val_1;
  assign DaRAT_val_2 = _zz_DaRAT_val_2;
  assign DaRAT_val_3 = _zz_DaRAT_val_3;
  assign DaRAT_val_4 = _zz_DaRAT_val_4;
  assign DaRAT_val_5 = _zz_DaRAT_val_5;
  assign DaRAT_val_6 = _zz_DaRAT_val_6;
  assign DaRAT_val_7 = _zz_DaRAT_val_7;
  assign DaRAT_val_8 = _zz_DaRAT_val_8;
  assign DaRAT_val_9 = _zz_DaRAT_val_9;
  assign DaRAT_val_10 = _zz_DaRAT_val_10;
  assign DaRAT_val_11 = _zz_DaRAT_val_11;
  assign DaRAT_val_12 = _zz_DaRAT_val_12;
  assign DaRAT_val_13 = _zz_DaRAT_val_13;
  assign DaRAT_val_14 = _zz_DaRAT_val_14;
  assign DaRAT_val_15 = _zz_DaRAT_val_15;
  assign DaRAT_val_16 = _zz_DaRAT_val_16;
  assign DaRAT_val_17 = _zz_DaRAT_val_17;
  assign DaRAT_val_18 = _zz_DaRAT_val_18;
  assign DaRAT_val_19 = _zz_DaRAT_val_19;
  assign DaRAT_val_20 = _zz_DaRAT_val_20;
  assign DaRAT_val_21 = _zz_DaRAT_val_21;
  assign DaRAT_val_22 = _zz_DaRAT_val_22;
  assign DaRAT_val_23 = _zz_DaRAT_val_23;
  assign DaRAT_val_24 = _zz_DaRAT_val_24;
  assign DaRAT_val_25 = _zz_DaRAT_val_25;
  assign DaRAT_val_26 = _zz_DaRAT_val_26;
  assign DaRAT_val_27 = _zz_DaRAT_val_27;
  assign DaRAT_val_28 = _zz_DaRAT_val_28;
  assign DaRAT_val_29 = _zz_DaRAT_val_29;
  assign DaRAT_val_30 = _zz_DaRAT_val_30;
  assign DaRAT_val_31 = _zz_DaRAT_val_31;
  assign DaRAT_val_0 = 32'h00000000;
  assign DifftestBundle_DifftestInstrCommitIndex_0 = 8'h00;
  assign DifftestBundle_DifftestInstrCommitIndex_1 = 8'h01;
  assign DifftestBundle_DifftestInstrCommitIndex_2 = 8'h02;
  assign DifftestBundle_DifftestInstrCommitIndex_3 = 8'h03;
  assign DifftestBundle_DifftestInstrCommitIndex_4 = 8'h04;
  assign DifftestBundle_DifftestInstrCommitValid_0 = cpuClockingArea_areaFlushReset_commitALU0_io_rob_valid;
  assign DifftestBundle_DifftestInstrCommitValid_1 = cpuClockingArea_areaFlushReset_commitALU1_io_rob_valid;
  assign DifftestBundle_DifftestInstrCommitValid_2 = cpuClockingArea_areaFlushReset_commitMULU_io_rob_valid;
  assign DifftestBundle_DifftestInstrCommitValid_3 = cpuClockingArea_areaFlushReset_commitDIVU_io_rob_valid;
  assign DifftestBundle_DifftestInstrCommitValid_4 = cpuClockingArea_areaFlushReset_commitLSU_io_rob_valid;
  assign DifftestBundle_DifftestInstrCommitPC_0 = {32'd0, _zz_DifftestBundle_DifftestInstrCommitPC_0};
  assign DifftestBundle_DifftestInstrCommitPC_1 = {32'd0, _zz_DifftestBundle_DifftestInstrCommitPC_1};
  assign DifftestBundle_DifftestInstrCommitPC_2 = {32'd0, _zz_DifftestBundle_DifftestInstrCommitPC_2};
  assign DifftestBundle_DifftestInstrCommitPC_3 = {32'd0, _zz_DifftestBundle_DifftestInstrCommitPC_3};
  assign DifftestBundle_DifftestInstrCommitPC_4 = {32'd0, _zz_DifftestBundle_DifftestInstrCommitPC_4};
  assign DifftestBundle_DifftestInstrCommitInstr_0 = 32'h00000000;
  assign DifftestBundle_DifftestInstrCommitInstr_1 = 32'h00000000;
  assign DifftestBundle_DifftestInstrCommitInstr_2 = 32'h00000000;
  assign DifftestBundle_DifftestInstrCommitInstr_3 = 32'h00000000;
  assign DifftestBundle_DifftestInstrCommitInstr_4 = 32'h00000000;
  assign DifftestBundle_DifftestSkip_0 = 1'b0;
  assign DifftestBundle_DifftestSkip_1 = 1'b0;
  assign DifftestBundle_DifftestSkip_2 = 1'b0;
  assign DifftestBundle_DifftestSkip_3 = 1'b0;
  assign DifftestBundle_DifftestSkip_4 = 1'b0;
  assign DifftestBundle_DifftestIsTlbFill_4 = (cpuClockingArea_memService_io_TLBCtrl_op == TLBOp_fill);
  assign DifftestBundle_DifftestTlbFillIndex_4 = {3'd0, _zz_DifftestBundle_DifftestTlbFillIndex_4};
  assign DifftestBundle_DifftestIsTlbFill_0 = 1'b0;
  assign DifftestBundle_DifftestTlbFillIndex_0 = 5'h00;
  assign DifftestBundle_DifftestIsTlbFill_1 = 1'b0;
  assign DifftestBundle_DifftestTlbFillIndex_1 = 5'h00;
  assign DifftestBundle_DifftestIsTlbFill_2 = 1'b0;
  assign DifftestBundle_DifftestTlbFillIndex_2 = 5'h00;
  assign DifftestBundle_DifftestIsTlbFill_3 = 1'b0;
  assign DifftestBundle_DifftestTlbFillIndex_3 = 5'h00;
  assign DifftestBundle_DifftestIsCount_1 = (cpuClockingArea_rob_io_commitROBEntries_1_specialOp == ROBSpecialOp_readCNT);
  assign DifftestBundle_DifftestCount_1 = {32'd0, _zz_DifftestBundle_DifftestCount_1};
  assign DifftestBundle_DifftestIsCount_2 = 1'b0;
  assign DifftestBundle_DifftestCount_2 = 64'h0000000000000000;
  assign DifftestBundle_DifftestIsCount_3 = 1'b0;
  assign DifftestBundle_DifftestCount_3 = 64'h0000000000000000;
  assign DifftestBundle_DifftestIsCount_4 = 1'b0;
  assign DifftestBundle_DifftestCount_4 = 64'h0000000000000000;
  assign DifftestBundle_DifftestIsCount_0 = 1'b0;
  assign DifftestBundle_DifftestCount_0 = 64'h0000000000000000;
  assign DifftestBundle_DifftestWen_0 = toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_valid;
  assign DifftestBundle_DifftestWen_1 = toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_valid;
  assign DifftestBundle_DifftestWen_2 = toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_valid;
  assign DifftestBundle_DifftestWen_3 = toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_valid;
  assign DifftestBundle_DifftestWen_4 = toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_valid;
  assign DifftestBundle_DifftestWdata_0 = {32'd0, _zz_DifftestBundle_DifftestWdata_0};
  assign DifftestBundle_DifftestWdata_1 = {32'd0, _zz_DifftestBundle_DifftestWdata_1};
  assign DifftestBundle_DifftestWdata_2 = {32'd0, _zz_DifftestBundle_DifftestWdata_2};
  assign DifftestBundle_DifftestWdata_3 = {32'd0, _zz_DifftestBundle_DifftestWdata_3};
  assign DifftestBundle_DifftestWdata_4 = {32'd0, _zz_DifftestBundle_DifftestWdata_4};
  assign DifftestBundle_DifftestWdest_0 = {2'd0, toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_m2sPipe_payload_prd};
  assign DifftestBundle_DifftestWdest_1 = {2'd0, toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_m2sPipe_payload_prd};
  assign DifftestBundle_DifftestWdest_2 = {2'd0, toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_m2sPipe_payload_prd};
  assign DifftestBundle_DifftestWdest_3 = {2'd0, toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_m2sPipe_payload_prd};
  assign DifftestBundle_DifftestWdest_4 = {2'd0, toplevel_cpuClockingArea_fuLSU_io_output_m2sPipe_payload_prd};
  assign DifftestBundle_DifftestCsrRstat_0 = ((cpuClockingArea_rob_io_commitROBEntries_0_specialOp == ROBSpecialOp_writeCSR) || (cpuClockingArea_rob_io_commitROBEntries_0_specialOp == ROBSpecialOp_readCSR));
  assign DifftestBundle_DifftestCsrData_0 = cpuClockingArea_csr_io_swRead_value;
  assign DifftestBundle_DifftestCsrRstat_1 = 1'b0;
  assign DifftestBundle_DifftestCsrData_1 = 32'h00000000;
  assign DifftestBundle_DifftestCsrRstat_2 = 1'b0;
  assign DifftestBundle_DifftestCsrData_2 = 32'h00000000;
  assign DifftestBundle_DifftestCsrRstat_3 = 1'b0;
  assign DifftestBundle_DifftestCsrData_3 = 32'h00000000;
  assign DifftestBundle_DifftestCsrRstat_4 = 1'b0;
  assign DifftestBundle_DifftestCsrData_4 = 32'h00000000;
  assign DifftestBundle_DifftestExcpEventExcpValid = (cpuClockingArea_rob_io_csrCtrl_tlbrException || cpuClockingArea_rob_io_csrCtrl_tlbrException);
  assign DifftestBundle_DifftestExcpEventEret = cpuClockingArea_rob_io_csrCtrl_ertn;
  assign DifftestBundle_DifftestExcpEventIntrNO = {24'd0, intrpt};
  assign DifftestBundle_DifftestExcpEventCause = {26'd0, cpuClockingArea_rob_io_csrCtrl_eCode};
  assign DifftestBundle_DifftestExcpEventEPC = {32'd0, _zz_DifftestBundle_DifftestExcpEventEPC};
  assign DifftestBundle_DifftestExcpEventInst = 32'h00000000;
  assign DifftestBundle_DifftestStoreEventData = {32'd0, cpuClockingArea_fuLSU_io_storeData};
  assign DifftestBundle_DifftestStoreEventValid = {4'd0, cpuClockingArea_fuLSU_io_storeMask};
  assign DifftestBundle_DifftestStoreEventVAddr = {32'd0, cpuClockingArea_fuLSU_io_VAddr};
  assign DifftestBundle_DifftestStoreEventPAddr = {32'd0, cpuClockingArea_fuLSU_io_PAddr};
  assign DifftestBundle_DifftestLoadEventValid = {4'd0, cpuClockingArea_fuLSU_io_loadMask};
  assign DifftestBundle_DifftestLoadEventVAddr = {32'd0, cpuClockingArea_fuLSU_io_VAddr};
  assign DifftestBundle_DifftestLoadEventPAddr = {32'd0, cpuClockingArea_fuLSU_io_PAddr};
  assign DifftestBundle_DifftestCSRRegStateCRMD = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_crmd};
  assign DifftestBundle_DifftestCSRRegStatePRMD = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_prmd};
  assign DifftestBundle_DifftestCSRRegStateECFG = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_ecfg};
  assign DifftestBundle_DifftestCSRRegStateESTAT = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_estat};
  assign DifftestBundle_DifftestCSRRegStateERA = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_era};
  assign DifftestBundle_DifftestCSRRegStateBADV = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_badv};
  assign DifftestBundle_DifftestCSRRegStateEENTRY = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_eentry};
  assign DifftestBundle_DifftestCSRRegStateTLBIDX = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_tlbidx};
  assign DifftestBundle_DifftestCSRRegStateTLBEHI = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_tlbehi};
  assign DifftestBundle_DifftestCSRRegStateTLBELO0 = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_tlbelo0};
  assign DifftestBundle_DifftestCSRRegStateTLBELO1 = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_tlbelo1};
  assign DifftestBundle_DifftestCSRRegStateASID = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_asid};
  assign DifftestBundle_DifftestCSRRegStatePGDL = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_pgdl};
  assign DifftestBundle_DifftestCSRRegStatePGDH = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_pgdh};
  assign DifftestBundle_DifftestCSRRegStateSAVE0 = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_save0};
  assign DifftestBundle_DifftestCSRRegStateSAVE1 = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_save1};
  assign DifftestBundle_DifftestCSRRegStateSAVE2 = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_save2};
  assign DifftestBundle_DifftestCSRRegStateSAVE3 = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_save3};
  assign DifftestBundle_DifftestCSRRegStateTID = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_tid};
  assign DifftestBundle_DifftestCSRRegStateTCFG = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_tcfg};
  assign DifftestBundle_DifftestCSRRegStateTVAL = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_tval};
  assign DifftestBundle_DifftestCSRRegStateTICLR = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_ticlr};
  assign DifftestBundle_DifftestCSRRegStateLLBCTL = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_llbctl};
  assign DifftestBundle_DifftestCSRRegStateTLBRENTRY = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_tlbrentry};
  assign DifftestBundle_DifftestCSRRegStateDMW0 = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_dmw0};
  assign DifftestBundle_DifftestCSRRegStateDMW1 = {32'd0, cpuClockingArea_csr_io_diffCSRBundle_dmw1};
  assign DifftestDelayBundle_DifftestInstrCommitIndex_0 = _zz_DifftestDelayBundle_DifftestInstrCommitIndex_0_1;
  assign DifftestDelayBundle_DifftestInstrCommitIndex_1 = _zz_DifftestDelayBundle_DifftestInstrCommitIndex_1_1;
  assign DifftestDelayBundle_DifftestInstrCommitIndex_2 = _zz_DifftestDelayBundle_DifftestInstrCommitIndex_2_1;
  assign DifftestDelayBundle_DifftestInstrCommitIndex_3 = _zz_DifftestDelayBundle_DifftestInstrCommitIndex_3_1;
  assign DifftestDelayBundle_DifftestInstrCommitIndex_4 = _zz_DifftestDelayBundle_DifftestInstrCommitIndex_4_1;
  assign DifftestDelayBundle_DifftestInstrCommitValid_0 = _zz_DifftestDelayBundle_DifftestInstrCommitValid_0_1;
  assign DifftestDelayBundle_DifftestInstrCommitValid_1 = _zz_DifftestDelayBundle_DifftestInstrCommitValid_1_1;
  assign DifftestDelayBundle_DifftestInstrCommitValid_2 = _zz_DifftestDelayBundle_DifftestInstrCommitValid_2_1;
  assign DifftestDelayBundle_DifftestInstrCommitValid_3 = _zz_DifftestDelayBundle_DifftestInstrCommitValid_3_1;
  assign DifftestDelayBundle_DifftestInstrCommitValid_4 = _zz_DifftestDelayBundle_DifftestInstrCommitValid_4_1;
  assign DifftestDelayBundle_DifftestInstrCommitPC_0 = _zz_DifftestDelayBundle_DifftestInstrCommitPC_0_1;
  assign DifftestDelayBundle_DifftestInstrCommitPC_1 = _zz_DifftestDelayBundle_DifftestInstrCommitPC_1_1;
  assign DifftestDelayBundle_DifftestInstrCommitPC_2 = _zz_DifftestDelayBundle_DifftestInstrCommitPC_2_1;
  assign DifftestDelayBundle_DifftestInstrCommitPC_3 = _zz_DifftestDelayBundle_DifftestInstrCommitPC_3_1;
  assign DifftestDelayBundle_DifftestInstrCommitPC_4 = _zz_DifftestDelayBundle_DifftestInstrCommitPC_4_1;
  assign DifftestDelayBundle_DifftestInstrCommitInstr_0 = _zz_DifftestDelayBundle_DifftestInstrCommitInstr_0_1;
  assign DifftestDelayBundle_DifftestInstrCommitInstr_1 = _zz_DifftestDelayBundle_DifftestInstrCommitInstr_1_1;
  assign DifftestDelayBundle_DifftestInstrCommitInstr_2 = _zz_DifftestDelayBundle_DifftestInstrCommitInstr_2_1;
  assign DifftestDelayBundle_DifftestInstrCommitInstr_3 = _zz_DifftestDelayBundle_DifftestInstrCommitInstr_3_1;
  assign DifftestDelayBundle_DifftestInstrCommitInstr_4 = _zz_DifftestDelayBundle_DifftestInstrCommitInstr_4_1;
  assign DifftestDelayBundle_DifftestSkip_0 = _zz_DifftestDelayBundle_DifftestSkip_0_1;
  assign DifftestDelayBundle_DifftestSkip_1 = _zz_DifftestDelayBundle_DifftestSkip_1_1;
  assign DifftestDelayBundle_DifftestSkip_2 = _zz_DifftestDelayBundle_DifftestSkip_2_1;
  assign DifftestDelayBundle_DifftestSkip_3 = _zz_DifftestDelayBundle_DifftestSkip_3_1;
  assign DifftestDelayBundle_DifftestSkip_4 = _zz_DifftestDelayBundle_DifftestSkip_4_1;
  assign DifftestDelayBundle_DifftestIsTlbFill_0 = _zz_DifftestDelayBundle_DifftestIsTlbFill_0_1;
  assign DifftestDelayBundle_DifftestIsTlbFill_1 = _zz_DifftestDelayBundle_DifftestIsTlbFill_1_1;
  assign DifftestDelayBundle_DifftestIsTlbFill_2 = _zz_DifftestDelayBundle_DifftestIsTlbFill_2_1;
  assign DifftestDelayBundle_DifftestIsTlbFill_3 = _zz_DifftestDelayBundle_DifftestIsTlbFill_3_1;
  assign DifftestDelayBundle_DifftestIsTlbFill_4 = _zz_DifftestDelayBundle_DifftestIsTlbFill_4_1;
  assign DifftestDelayBundle_DifftestTlbFillIndex_0 = _zz_DifftestDelayBundle_DifftestTlbFillIndex_0_1;
  assign DifftestDelayBundle_DifftestTlbFillIndex_1 = _zz_DifftestDelayBundle_DifftestTlbFillIndex_1_1;
  assign DifftestDelayBundle_DifftestTlbFillIndex_2 = _zz_DifftestDelayBundle_DifftestTlbFillIndex_2_1;
  assign DifftestDelayBundle_DifftestTlbFillIndex_3 = _zz_DifftestDelayBundle_DifftestTlbFillIndex_3_1;
  assign DifftestDelayBundle_DifftestTlbFillIndex_4 = _zz_DifftestDelayBundle_DifftestTlbFillIndex_4_1;
  assign DifftestDelayBundle_DifftestIsCount_0 = _zz_DifftestDelayBundle_DifftestIsCount_0_1;
  assign DifftestDelayBundle_DifftestIsCount_1 = _zz_DifftestDelayBundle_DifftestIsCount_1_1;
  assign DifftestDelayBundle_DifftestIsCount_2 = _zz_DifftestDelayBundle_DifftestIsCount_2_1;
  assign DifftestDelayBundle_DifftestIsCount_3 = _zz_DifftestDelayBundle_DifftestIsCount_3_1;
  assign DifftestDelayBundle_DifftestIsCount_4 = _zz_DifftestDelayBundle_DifftestIsCount_4_1;
  assign DifftestDelayBundle_DifftestCount_0 = _zz_DifftestDelayBundle_DifftestCount_0_1;
  assign DifftestDelayBundle_DifftestCount_1 = _zz_DifftestDelayBundle_DifftestCount_1_1;
  assign DifftestDelayBundle_DifftestCount_2 = _zz_DifftestDelayBundle_DifftestCount_2_1;
  assign DifftestDelayBundle_DifftestCount_3 = _zz_DifftestDelayBundle_DifftestCount_3_1;
  assign DifftestDelayBundle_DifftestCount_4 = _zz_DifftestDelayBundle_DifftestCount_4_1;
  assign DifftestDelayBundle_DifftestWen_0 = _zz_DifftestDelayBundle_DifftestWen_0_1;
  assign DifftestDelayBundle_DifftestWen_1 = _zz_DifftestDelayBundle_DifftestWen_1_1;
  assign DifftestDelayBundle_DifftestWen_2 = _zz_DifftestDelayBundle_DifftestWen_2_1;
  assign DifftestDelayBundle_DifftestWen_3 = _zz_DifftestDelayBundle_DifftestWen_3_1;
  assign DifftestDelayBundle_DifftestWen_4 = _zz_DifftestDelayBundle_DifftestWen_4_1;
  assign DifftestDelayBundle_DifftestWdest_0 = _zz_DifftestDelayBundle_DifftestWdest_0_1;
  assign DifftestDelayBundle_DifftestWdest_1 = _zz_DifftestDelayBundle_DifftestWdest_1_1;
  assign DifftestDelayBundle_DifftestWdest_2 = _zz_DifftestDelayBundle_DifftestWdest_2_1;
  assign DifftestDelayBundle_DifftestWdest_3 = _zz_DifftestDelayBundle_DifftestWdest_3_1;
  assign DifftestDelayBundle_DifftestWdest_4 = _zz_DifftestDelayBundle_DifftestWdest_4_1;
  assign DifftestDelayBundle_DifftestWdata_0 = _zz_DifftestDelayBundle_DifftestWdata_0_1;
  assign DifftestDelayBundle_DifftestWdata_1 = _zz_DifftestDelayBundle_DifftestWdata_1_1;
  assign DifftestDelayBundle_DifftestWdata_2 = _zz_DifftestDelayBundle_DifftestWdata_2_1;
  assign DifftestDelayBundle_DifftestWdata_3 = _zz_DifftestDelayBundle_DifftestWdata_3_1;
  assign DifftestDelayBundle_DifftestWdata_4 = _zz_DifftestDelayBundle_DifftestWdata_4_1;
  assign DifftestDelayBundle_DifftestCsrRstat_0 = _zz_DifftestDelayBundle_DifftestCsrRstat_0_1;
  assign DifftestDelayBundle_DifftestCsrRstat_1 = _zz_DifftestDelayBundle_DifftestCsrRstat_1_1;
  assign DifftestDelayBundle_DifftestCsrRstat_2 = _zz_DifftestDelayBundle_DifftestCsrRstat_2_1;
  assign DifftestDelayBundle_DifftestCsrRstat_3 = _zz_DifftestDelayBundle_DifftestCsrRstat_3_1;
  assign DifftestDelayBundle_DifftestCsrRstat_4 = _zz_DifftestDelayBundle_DifftestCsrRstat_4_1;
  assign DifftestDelayBundle_DifftestCsrData_0 = _zz_DifftestDelayBundle_DifftestCsrData_0_1;
  assign DifftestDelayBundle_DifftestCsrData_1 = _zz_DifftestDelayBundle_DifftestCsrData_1_1;
  assign DifftestDelayBundle_DifftestCsrData_2 = _zz_DifftestDelayBundle_DifftestCsrData_2_1;
  assign DifftestDelayBundle_DifftestCsrData_3 = _zz_DifftestDelayBundle_DifftestCsrData_3_1;
  assign DifftestDelayBundle_DifftestCsrData_4 = _zz_DifftestDelayBundle_DifftestCsrData_4_1;
  assign DifftestDelayBundle_DifftestExcpEventExcpValid = _zz_DifftestDelayBundle_DifftestExcpEventExcpValid_1;
  assign DifftestDelayBundle_DifftestExcpEventEret = _zz_DifftestDelayBundle_DifftestExcpEventEret_1;
  assign DifftestDelayBundle_DifftestExcpEventIntrNO = _zz_DifftestDelayBundle_DifftestExcpEventIntrNO_1;
  assign DifftestDelayBundle_DifftestExcpEventCause = _zz_DifftestDelayBundle_DifftestExcpEventCause_1;
  assign DifftestDelayBundle_DifftestExcpEventEPC = _zz_DifftestDelayBundle_DifftestExcpEventEPC_1;
  assign DifftestDelayBundle_DifftestExcpEventInst = _zz_DifftestDelayBundle_DifftestExcpEventInst_1;
  assign DifftestDelayBundle_DifftestStoreEventValid = _zz_DifftestDelayBundle_DifftestStoreEventValid_1;
  assign DifftestDelayBundle_DifftestStoreEventPAddr = _zz_DifftestDelayBundle_DifftestStoreEventPAddr_1;
  assign DifftestDelayBundle_DifftestStoreEventVAddr = _zz_DifftestDelayBundle_DifftestStoreEventVAddr_1;
  assign DifftestDelayBundle_DifftestStoreEventData = _zz_DifftestDelayBundle_DifftestStoreEventData_1;
  assign DifftestDelayBundle_DifftestLoadEventValid = _zz_DifftestDelayBundle_DifftestLoadEventValid_1;
  assign DifftestDelayBundle_DifftestLoadEventPAddr = _zz_DifftestDelayBundle_DifftestLoadEventPAddr_1;
  assign DifftestDelayBundle_DifftestLoadEventVAddr = _zz_DifftestDelayBundle_DifftestLoadEventVAddr_1;
  assign arid = cpuClockingArea_arbiter_io_out_arid;
  assign araddr = cpuClockingArea_arbiter_io_out_araddr;
  assign arlen = cpuClockingArea_arbiter_io_out_arlen;
  assign arsize = cpuClockingArea_arbiter_io_out_arsize;
  assign arburst = cpuClockingArea_arbiter_io_out_arburst;
  assign arlock = cpuClockingArea_arbiter_io_out_arlock;
  assign arcache = cpuClockingArea_arbiter_io_out_arcache;
  assign arprot = cpuClockingArea_arbiter_io_out_arprot;
  assign arvalid = cpuClockingArea_arbiter_io_out_arvalid;
  assign rready = cpuClockingArea_arbiter_io_out_rready;
  assign awid = cpuClockingArea_arbiter_io_out_awid;
  assign awaddr = cpuClockingArea_arbiter_io_out_awaddr;
  assign awlen = cpuClockingArea_arbiter_io_out_awlen;
  assign awsize = cpuClockingArea_arbiter_io_out_awsize;
  assign awburst = cpuClockingArea_arbiter_io_out_awburst;
  assign awlock = cpuClockingArea_arbiter_io_out_awlock;
  assign awcache = cpuClockingArea_arbiter_io_out_awcache;
  assign awprot = cpuClockingArea_arbiter_io_out_awprot;
  assign awvalid = cpuClockingArea_arbiter_io_out_awvalid;
  assign wid = cpuClockingArea_arbiter_io_out_wid;
  assign wdata = cpuClockingArea_arbiter_io_out_wdata;
  assign wstrb = cpuClockingArea_arbiter_io_out_wstrb;
  assign wlast = cpuClockingArea_arbiter_io_out_wlast;
  assign wvalid = cpuClockingArea_arbiter_io_out_wvalid;
  assign bready = cpuClockingArea_arbiter_io_out_bready;
  assign debug0_wb_pc = 32'h00000000;
  assign debug0_wb_rf_wen = 4'b0000;
  assign debug0_wb_rf_wnum = 5'h00;
  assign debug0_wb_rf_wdata = 32'h00000000;
  assign ws_valid = 1'b0;
  assign rf_rdata = 32'h00000000;
  always @(posedge aclk) begin
    if(!cpuClockingArea_areaFlushReset_newReset) begin
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rValid <= 1'b0;
      toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rValid <= 1'b0;
      toplevel_cpuClockingArea_fuLSU_io_output_rValid <= 1'b0;
    end else begin
      if(cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rValid <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_valid;
      end
      if(cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rValid <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_valid;
      end
      if(cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rValid <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_valid;
      end
      if(cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rValid <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_valid;
      end
      if(cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rValid <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_valid;
      end
      if(cpuClockingArea_areaFlushReset_roALU0_io_toFU_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rValid <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_valid;
      end
      if(cpuClockingArea_areaFlushReset_roALU1_io_toFU_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rValid <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_valid;
      end
      if(cpuClockingArea_areaFlushReset_roMULU_io_toFU_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rValid <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_valid;
      end
      if(cpuClockingArea_areaFlushReset_roDIVU_io_toFU_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rValid <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_valid;
      end
      if(cpuClockingArea_areaFlushReset_roLSU_io_toFU_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rValid <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_valid;
      end
      if(cpuClockingArea_areaFlushReset_fuALU0_io_output_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rValid <= cpuClockingArea_areaFlushReset_fuALU0_io_output_valid;
      end
      if(cpuClockingArea_areaFlushReset_fuALU1_io_output_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rValid <= cpuClockingArea_areaFlushReset_fuALU1_io_output_valid;
      end
      if(cpuClockingArea_areaFlushReset_fuMULU_io_output_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rValid <= cpuClockingArea_areaFlushReset_fuMULU_io_output_valid;
      end
      if(cpuClockingArea_areaFlushReset_fuDIVU_io_output_ready) begin
        toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rValid <= cpuClockingArea_areaFlushReset_fuDIVU_io_output_valid;
      end
      if(cpuClockingArea_fuLSU_io_output_ready) begin
        toplevel_cpuClockingArea_fuLSU_io_output_rValid <= cpuClockingArea_fuLSU_io_output_valid;
      end
    end
  end

  always @(posedge aclk) begin
    if(cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_robIdx <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_branchInfo_predictPC <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_branchInfo_predictPC;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_branchInfo_predictResult <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_branchInfo_predictResult;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_exceptionInfo_eSubCode;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_pc <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_pc;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_prd <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_psrc_0 <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_psrc_0;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_psrc_1 <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_psrc_1;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_imm <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_imm;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_aluOp <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_uop_aluOp;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_bruOp <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_uop_bruOp;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_uop_cruOp <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_uop_cruOp;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_rData_roop_aluROOp <= cpuClockingArea_areaFlushReset_issueQueueALU0_io_output_payload_roop_aluROOp;
    end
    if(cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_robIdx <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_branchInfo_predictPC <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_branchInfo_predictPC;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_branchInfo_predictResult <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_branchInfo_predictResult;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_exceptionInfo_eSubCode;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_pc <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_pc;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_prd <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_psrc_0 <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_psrc_0;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_psrc_1 <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_psrc_1;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_imm <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_imm;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_aluOp <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_uop_aluOp;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_uop_bruOp <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_uop_bruOp;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_aluROOp <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_roop_aluROOp;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_rData_roop_cruROOp <= cpuClockingArea_areaFlushReset_issueQueueALU1_io_output_payload_roop_cruROOp;
    end
    if(cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_robIdx <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_branchResult_targetPC <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_branchResult_targetPC;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_branchResult_branchResult <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_branchResult_branchResult;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_branchResult_predictFail <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_branchResult_predictFail;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_exceptionInfo_eSubCode;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_pc <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_pc;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_prd <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_psrc_0 <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_psrc_0;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_psrc_1 <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_psrc_1;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_imm <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_imm;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_rData_uop_muluOp <= cpuClockingArea_areaFlushReset_issueQueueMULU_io_output_payload_uop_muluOp;
    end
    if(cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_robIdx <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_branchResult_targetPC <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_branchResult_targetPC;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_branchResult_branchResult <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_branchResult_branchResult;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_branchResult_predictFail <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_branchResult_predictFail;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_exceptionInfo_eSubCode;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_pc <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_pc;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_prd <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_psrc_0 <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_psrc_0;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_psrc_1 <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_psrc_1;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_imm <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_imm;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_rData_uop_divuOp <= cpuClockingArea_areaFlushReset_issueQueueDIVU_io_output_payload_uop_divuOp;
    end
    if(cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_robIdx <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_branchResult_targetPC <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_branchResult_targetPC;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_branchResult_branchResult <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_branchResult_branchResult;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_branchResult_predictFail <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_branchResult_predictFail;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_exceptionInfo_eSubCode;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_pc <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_pc;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_prd <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_psrc_0 <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_psrc_0;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_psrc_1 <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_psrc_1;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_imm <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_imm;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuOp <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_uop_lsuOp;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_uop_lsuCoOp <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_uop_lsuCoOp;
      toplevel_cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_rData_roop_lsuROOp <= cpuClockingArea_areaFlushReset_issueQueueLSU_io_output_payload_roop_lsuROOp;
    end
    if(cpuClockingArea_areaFlushReset_roALU0_io_toFU_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src1 <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src1;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src2 <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src2;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src3 <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src3;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_src4 <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_src4;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_robIdx <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_branchInfo_predictPC <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_branchInfo_predictPC;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_branchInfo_predictResult <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_branchInfo_predictResult;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_exceptionInfo_eSubCode;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_pc <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_pc;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_prd <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_aluOp <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_uop_aluOp;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_bruOp <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_uop_bruOp;
      toplevel_cpuClockingArea_areaFlushReset_roALU0_io_toFU_rData_uop_cruOp <= cpuClockingArea_areaFlushReset_roALU0_io_toFU_payload_uop_cruOp;
    end
    if(cpuClockingArea_areaFlushReset_roALU1_io_toFU_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src1 <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src1;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src2 <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src2;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src3 <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src3;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_src4 <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_src4;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_robIdx <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_branchInfo_predictPC <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_branchInfo_predictPC;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_branchInfo_predictResult <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_branchInfo_predictResult;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_exceptionInfo_eSubCode;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_pc <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_pc;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_prd <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_aluOp <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_uop_aluOp;
      toplevel_cpuClockingArea_areaFlushReset_roALU1_io_toFU_rData_uop_bruOp <= cpuClockingArea_areaFlushReset_roALU1_io_toFU_payload_uop_bruOp;
    end
    if(cpuClockingArea_areaFlushReset_roMULU_io_toFU_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_src1 <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_src1;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_src2 <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_src2;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_robIdx <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_branchResult_targetPC <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_branchResult_targetPC;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_branchResult_branchResult <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_branchResult_branchResult;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_branchResult_predictFail <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_branchResult_predictFail;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_exceptionInfo_eSubCode;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_pc <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_pc;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_prd <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_roMULU_io_toFU_rData_uop_muluOp <= cpuClockingArea_areaFlushReset_roMULU_io_toFU_payload_uop_muluOp;
    end
    if(cpuClockingArea_areaFlushReset_roDIVU_io_toFU_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_src1 <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_src1;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_src2 <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_src2;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_robIdx <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_branchResult_targetPC <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_branchResult_targetPC;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_branchResult_branchResult <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_branchResult_branchResult;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_branchResult_predictFail <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_branchResult_predictFail;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_exceptionInfo_eSubCode;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_pc <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_pc;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_prd <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_roDIVU_io_toFU_rData_uop_divuOp <= cpuClockingArea_areaFlushReset_roDIVU_io_toFU_payload_uop_divuOp;
    end
    if(cpuClockingArea_areaFlushReset_roLSU_io_toFU_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_src1 <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_src1;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_src2 <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_src2;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_src3 <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_src3;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_robIdx <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_branchResult_targetPC <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_branchResult_targetPC;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_branchResult_branchResult <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_branchResult_branchResult;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_branchResult_predictFail <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_branchResult_predictFail;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_exceptionInfo_eSubCode;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_pc <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_pc;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_prd <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuOp <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_uop_lsuOp;
      toplevel_cpuClockingArea_areaFlushReset_roLSU_io_toFU_rData_uop_lsuCoOp <= cpuClockingArea_areaFlushReset_roLSU_io_toFU_payload_uop_lsuCoOp;
    end
    if(cpuClockingArea_areaFlushReset_fuALU0_io_output_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_robIdx <= cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_data <= cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_data;
      toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_prd <= cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_branchResult_targetPC <= cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_branchResult_targetPC;
      toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_branchResult_branchResult <= cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_branchResult_branchResult;
      toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_branchResult_predictFail <= cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_branchResult_predictFail;
      toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_fuALU0_io_output_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_fuALU0_io_output_payload_exceptionInfo_eSubCode;
    end
    if(cpuClockingArea_areaFlushReset_fuALU1_io_output_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_robIdx <= cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_data <= cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_data;
      toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_prd <= cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_branchResult_targetPC <= cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_branchResult_targetPC;
      toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_branchResult_branchResult <= cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_branchResult_branchResult;
      toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_branchResult_predictFail <= cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_branchResult_predictFail;
      toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_fuALU1_io_output_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_fuALU1_io_output_payload_exceptionInfo_eSubCode;
    end
    if(cpuClockingArea_areaFlushReset_fuMULU_io_output_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_robIdx <= cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_data <= cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_data;
      toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_prd <= cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_branchResult_targetPC <= cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_branchResult_targetPC;
      toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_branchResult_branchResult <= cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_branchResult_branchResult;
      toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_branchResult_predictFail <= cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_branchResult_predictFail;
      toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_fuMULU_io_output_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_fuMULU_io_output_payload_exceptionInfo_eSubCode;
    end
    if(cpuClockingArea_areaFlushReset_fuDIVU_io_output_ready) begin
      toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_robIdx <= cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_robIdx;
      toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_data <= cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_data;
      toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_prd <= cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_prd;
      toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_branchResult_targetPC <= cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_branchResult_targetPC;
      toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_branchResult_branchResult <= cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_branchResult_branchResult;
      toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_branchResult_predictFail <= cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_branchResult_predictFail;
      toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_exceptionInfo_exception <= cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_exceptionInfo_eCode <= cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_areaFlushReset_fuDIVU_io_output_rData_exceptionInfo_eSubCode <= cpuClockingArea_areaFlushReset_fuDIVU_io_output_payload_exceptionInfo_eSubCode;
    end
    if(cpuClockingArea_fuLSU_io_output_ready) begin
      toplevel_cpuClockingArea_fuLSU_io_output_rData_robIdx <= cpuClockingArea_fuLSU_io_output_payload_robIdx;
      toplevel_cpuClockingArea_fuLSU_io_output_rData_data <= cpuClockingArea_fuLSU_io_output_payload_data;
      toplevel_cpuClockingArea_fuLSU_io_output_rData_prd <= cpuClockingArea_fuLSU_io_output_payload_prd;
      toplevel_cpuClockingArea_fuLSU_io_output_rData_branchResult_targetPC <= cpuClockingArea_fuLSU_io_output_payload_branchResult_targetPC;
      toplevel_cpuClockingArea_fuLSU_io_output_rData_branchResult_branchResult <= cpuClockingArea_fuLSU_io_output_payload_branchResult_branchResult;
      toplevel_cpuClockingArea_fuLSU_io_output_rData_branchResult_predictFail <= cpuClockingArea_fuLSU_io_output_payload_branchResult_predictFail;
      toplevel_cpuClockingArea_fuLSU_io_output_rData_exceptionInfo_exception <= cpuClockingArea_fuLSU_io_output_payload_exceptionInfo_exception;
      toplevel_cpuClockingArea_fuLSU_io_output_rData_exceptionInfo_eCode <= cpuClockingArea_fuLSU_io_output_payload_exceptionInfo_eCode;
      toplevel_cpuClockingArea_fuLSU_io_output_rData_exceptionInfo_eSubCode <= cpuClockingArea_fuLSU_io_output_payload_exceptionInfo_eSubCode;
    end
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_0 <= DifftestBundle_DifftestInstrCommitIndex_0;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_1 <= DifftestBundle_DifftestInstrCommitIndex_1;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_2 <= DifftestBundle_DifftestInstrCommitIndex_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_3 <= DifftestBundle_DifftestInstrCommitIndex_3;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_4 <= DifftestBundle_DifftestInstrCommitIndex_4;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_0 <= DifftestBundle_DifftestInstrCommitValid_0;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_1 <= DifftestBundle_DifftestInstrCommitValid_1;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_2 <= DifftestBundle_DifftestInstrCommitValid_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_3 <= DifftestBundle_DifftestInstrCommitValid_3;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_4 <= DifftestBundle_DifftestInstrCommitValid_4;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_0 <= DifftestBundle_DifftestInstrCommitPC_0;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_1 <= DifftestBundle_DifftestInstrCommitPC_1;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_2 <= DifftestBundle_DifftestInstrCommitPC_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_3 <= DifftestBundle_DifftestInstrCommitPC_3;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_4 <= DifftestBundle_DifftestInstrCommitPC_4;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_0 <= DifftestBundle_DifftestInstrCommitInstr_0;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_1 <= DifftestBundle_DifftestInstrCommitInstr_1;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_2 <= DifftestBundle_DifftestInstrCommitInstr_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_3 <= DifftestBundle_DifftestInstrCommitInstr_3;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_4 <= DifftestBundle_DifftestInstrCommitInstr_4;
    _zz_DifftestDelayBundle_DifftestSkip_0 <= DifftestBundle_DifftestSkip_0;
    _zz_DifftestDelayBundle_DifftestSkip_1 <= DifftestBundle_DifftestSkip_1;
    _zz_DifftestDelayBundle_DifftestSkip_2 <= DifftestBundle_DifftestSkip_2;
    _zz_DifftestDelayBundle_DifftestSkip_3 <= DifftestBundle_DifftestSkip_3;
    _zz_DifftestDelayBundle_DifftestSkip_4 <= DifftestBundle_DifftestSkip_4;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_0 <= DifftestBundle_DifftestIsTlbFill_0;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_1 <= DifftestBundle_DifftestIsTlbFill_1;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_2 <= DifftestBundle_DifftestIsTlbFill_2;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_3 <= DifftestBundle_DifftestIsTlbFill_3;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_4 <= DifftestBundle_DifftestIsTlbFill_4;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_0 <= DifftestBundle_DifftestTlbFillIndex_0;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_1 <= DifftestBundle_DifftestTlbFillIndex_1;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_2 <= DifftestBundle_DifftestTlbFillIndex_2;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_3 <= DifftestBundle_DifftestTlbFillIndex_3;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_4 <= DifftestBundle_DifftestTlbFillIndex_4;
    _zz_DifftestDelayBundle_DifftestIsCount_0 <= DifftestBundle_DifftestIsCount_0;
    _zz_DifftestDelayBundle_DifftestIsCount_1 <= DifftestBundle_DifftestIsCount_1;
    _zz_DifftestDelayBundle_DifftestIsCount_2 <= DifftestBundle_DifftestIsCount_2;
    _zz_DifftestDelayBundle_DifftestIsCount_3 <= DifftestBundle_DifftestIsCount_3;
    _zz_DifftestDelayBundle_DifftestIsCount_4 <= DifftestBundle_DifftestIsCount_4;
    _zz_DifftestDelayBundle_DifftestCount_0 <= DifftestBundle_DifftestCount_0;
    _zz_DifftestDelayBundle_DifftestCount_1 <= DifftestBundle_DifftestCount_1;
    _zz_DifftestDelayBundle_DifftestCount_2 <= DifftestBundle_DifftestCount_2;
    _zz_DifftestDelayBundle_DifftestCount_3 <= DifftestBundle_DifftestCount_3;
    _zz_DifftestDelayBundle_DifftestCount_4 <= DifftestBundle_DifftestCount_4;
    _zz_DifftestDelayBundle_DifftestWen_0 <= DifftestBundle_DifftestWen_0;
    _zz_DifftestDelayBundle_DifftestWen_1 <= DifftestBundle_DifftestWen_1;
    _zz_DifftestDelayBundle_DifftestWen_2 <= DifftestBundle_DifftestWen_2;
    _zz_DifftestDelayBundle_DifftestWen_3 <= DifftestBundle_DifftestWen_3;
    _zz_DifftestDelayBundle_DifftestWen_4 <= DifftestBundle_DifftestWen_4;
    _zz_DifftestDelayBundle_DifftestWdest_0 <= DifftestBundle_DifftestWdest_0;
    _zz_DifftestDelayBundle_DifftestWdest_1 <= DifftestBundle_DifftestWdest_1;
    _zz_DifftestDelayBundle_DifftestWdest_2 <= DifftestBundle_DifftestWdest_2;
    _zz_DifftestDelayBundle_DifftestWdest_3 <= DifftestBundle_DifftestWdest_3;
    _zz_DifftestDelayBundle_DifftestWdest_4 <= DifftestBundle_DifftestWdest_4;
    _zz_DifftestDelayBundle_DifftestWdata_0 <= DifftestBundle_DifftestWdata_0;
    _zz_DifftestDelayBundle_DifftestWdata_1 <= DifftestBundle_DifftestWdata_1;
    _zz_DifftestDelayBundle_DifftestWdata_2 <= DifftestBundle_DifftestWdata_2;
    _zz_DifftestDelayBundle_DifftestWdata_3 <= DifftestBundle_DifftestWdata_3;
    _zz_DifftestDelayBundle_DifftestWdata_4 <= DifftestBundle_DifftestWdata_4;
    _zz_DifftestDelayBundle_DifftestCsrRstat_0 <= DifftestBundle_DifftestCsrRstat_0;
    _zz_DifftestDelayBundle_DifftestCsrRstat_1 <= DifftestBundle_DifftestCsrRstat_1;
    _zz_DifftestDelayBundle_DifftestCsrRstat_2 <= DifftestBundle_DifftestCsrRstat_2;
    _zz_DifftestDelayBundle_DifftestCsrRstat_3 <= DifftestBundle_DifftestCsrRstat_3;
    _zz_DifftestDelayBundle_DifftestCsrRstat_4 <= DifftestBundle_DifftestCsrRstat_4;
    _zz_DifftestDelayBundle_DifftestCsrData_0 <= DifftestBundle_DifftestCsrData_0;
    _zz_DifftestDelayBundle_DifftestCsrData_1 <= DifftestBundle_DifftestCsrData_1;
    _zz_DifftestDelayBundle_DifftestCsrData_2 <= DifftestBundle_DifftestCsrData_2;
    _zz_DifftestDelayBundle_DifftestCsrData_3 <= DifftestBundle_DifftestCsrData_3;
    _zz_DifftestDelayBundle_DifftestCsrData_4 <= DifftestBundle_DifftestCsrData_4;
    _zz_DifftestDelayBundle_DifftestExcpEventExcpValid <= DifftestBundle_DifftestExcpEventExcpValid;
    _zz_DifftestDelayBundle_DifftestExcpEventEret <= DifftestBundle_DifftestExcpEventEret;
    _zz_DifftestDelayBundle_DifftestExcpEventIntrNO <= DifftestBundle_DifftestExcpEventIntrNO;
    _zz_DifftestDelayBundle_DifftestExcpEventCause <= DifftestBundle_DifftestExcpEventCause;
    _zz_DifftestDelayBundle_DifftestExcpEventEPC <= DifftestBundle_DifftestExcpEventEPC;
    _zz_DifftestDelayBundle_DifftestExcpEventInst <= DifftestBundle_DifftestExcpEventInst;
    _zz_DifftestDelayBundle_DifftestStoreEventValid <= DifftestBundle_DifftestStoreEventValid;
    _zz_DifftestDelayBundle_DifftestStoreEventPAddr <= DifftestBundle_DifftestStoreEventPAddr;
    _zz_DifftestDelayBundle_DifftestStoreEventVAddr <= DifftestBundle_DifftestStoreEventVAddr;
    _zz_DifftestDelayBundle_DifftestStoreEventData <= DifftestBundle_DifftestStoreEventData;
    _zz_DifftestDelayBundle_DifftestLoadEventValid <= DifftestBundle_DifftestLoadEventValid;
    _zz_DifftestDelayBundle_DifftestLoadEventPAddr <= DifftestBundle_DifftestLoadEventPAddr;
    _zz_DifftestDelayBundle_DifftestLoadEventVAddr <= DifftestBundle_DifftestLoadEventVAddr;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_0_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitIndex_0;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_1_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitIndex_1;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_2_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitIndex_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_3_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitIndex_3;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_4_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitIndex_4;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_0_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitValid_0;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_1_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitValid_1;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_2_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitValid_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_3_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitValid_3;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_4_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitValid_4;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_0_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitPC_0;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_1_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitPC_1;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_2_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitPC_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_3_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitPC_3;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_4_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitPC_4;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_0_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitInstr_0;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_1_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitInstr_1;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_2_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitInstr_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_3_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitInstr_3;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_4_2 <= _zz_DifftestDelayBundle_DifftestInstrCommitInstr_4;
    _zz_DifftestDelayBundle_DifftestSkip_0_2 <= _zz_DifftestDelayBundle_DifftestSkip_0;
    _zz_DifftestDelayBundle_DifftestSkip_1_2 <= _zz_DifftestDelayBundle_DifftestSkip_1;
    _zz_DifftestDelayBundle_DifftestSkip_2_2 <= _zz_DifftestDelayBundle_DifftestSkip_2;
    _zz_DifftestDelayBundle_DifftestSkip_3_2 <= _zz_DifftestDelayBundle_DifftestSkip_3;
    _zz_DifftestDelayBundle_DifftestSkip_4_2 <= _zz_DifftestDelayBundle_DifftestSkip_4;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_0_2 <= _zz_DifftestDelayBundle_DifftestIsTlbFill_0;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_1_2 <= _zz_DifftestDelayBundle_DifftestIsTlbFill_1;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_2_2 <= _zz_DifftestDelayBundle_DifftestIsTlbFill_2;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_3_2 <= _zz_DifftestDelayBundle_DifftestIsTlbFill_3;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_4_2 <= _zz_DifftestDelayBundle_DifftestIsTlbFill_4;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_0_2 <= _zz_DifftestDelayBundle_DifftestTlbFillIndex_0;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_1_2 <= _zz_DifftestDelayBundle_DifftestTlbFillIndex_1;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_2_2 <= _zz_DifftestDelayBundle_DifftestTlbFillIndex_2;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_3_2 <= _zz_DifftestDelayBundle_DifftestTlbFillIndex_3;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_4_2 <= _zz_DifftestDelayBundle_DifftestTlbFillIndex_4;
    _zz_DifftestDelayBundle_DifftestIsCount_0_2 <= _zz_DifftestDelayBundle_DifftestIsCount_0;
    _zz_DifftestDelayBundle_DifftestIsCount_1_2 <= _zz_DifftestDelayBundle_DifftestIsCount_1;
    _zz_DifftestDelayBundle_DifftestIsCount_2_2 <= _zz_DifftestDelayBundle_DifftestIsCount_2;
    _zz_DifftestDelayBundle_DifftestIsCount_3_2 <= _zz_DifftestDelayBundle_DifftestIsCount_3;
    _zz_DifftestDelayBundle_DifftestIsCount_4_2 <= _zz_DifftestDelayBundle_DifftestIsCount_4;
    _zz_DifftestDelayBundle_DifftestCount_0_2 <= _zz_DifftestDelayBundle_DifftestCount_0;
    _zz_DifftestDelayBundle_DifftestCount_1_2 <= _zz_DifftestDelayBundle_DifftestCount_1;
    _zz_DifftestDelayBundle_DifftestCount_2_2 <= _zz_DifftestDelayBundle_DifftestCount_2;
    _zz_DifftestDelayBundle_DifftestCount_3_2 <= _zz_DifftestDelayBundle_DifftestCount_3;
    _zz_DifftestDelayBundle_DifftestCount_4_2 <= _zz_DifftestDelayBundle_DifftestCount_4;
    _zz_DifftestDelayBundle_DifftestWen_0_2 <= _zz_DifftestDelayBundle_DifftestWen_0;
    _zz_DifftestDelayBundle_DifftestWen_1_2 <= _zz_DifftestDelayBundle_DifftestWen_1;
    _zz_DifftestDelayBundle_DifftestWen_2_2 <= _zz_DifftestDelayBundle_DifftestWen_2;
    _zz_DifftestDelayBundle_DifftestWen_3_2 <= _zz_DifftestDelayBundle_DifftestWen_3;
    _zz_DifftestDelayBundle_DifftestWen_4_2 <= _zz_DifftestDelayBundle_DifftestWen_4;
    _zz_DifftestDelayBundle_DifftestWdest_0_2 <= _zz_DifftestDelayBundle_DifftestWdest_0;
    _zz_DifftestDelayBundle_DifftestWdest_1_2 <= _zz_DifftestDelayBundle_DifftestWdest_1;
    _zz_DifftestDelayBundle_DifftestWdest_2_2 <= _zz_DifftestDelayBundle_DifftestWdest_2;
    _zz_DifftestDelayBundle_DifftestWdest_3_2 <= _zz_DifftestDelayBundle_DifftestWdest_3;
    _zz_DifftestDelayBundle_DifftestWdest_4_2 <= _zz_DifftestDelayBundle_DifftestWdest_4;
    _zz_DifftestDelayBundle_DifftestWdata_0_2 <= _zz_DifftestDelayBundle_DifftestWdata_0;
    _zz_DifftestDelayBundle_DifftestWdata_1_2 <= _zz_DifftestDelayBundle_DifftestWdata_1;
    _zz_DifftestDelayBundle_DifftestWdata_2_2 <= _zz_DifftestDelayBundle_DifftestWdata_2;
    _zz_DifftestDelayBundle_DifftestWdata_3_2 <= _zz_DifftestDelayBundle_DifftestWdata_3;
    _zz_DifftestDelayBundle_DifftestWdata_4_2 <= _zz_DifftestDelayBundle_DifftestWdata_4;
    _zz_DifftestDelayBundle_DifftestCsrRstat_0_2 <= _zz_DifftestDelayBundle_DifftestCsrRstat_0;
    _zz_DifftestDelayBundle_DifftestCsrRstat_1_2 <= _zz_DifftestDelayBundle_DifftestCsrRstat_1;
    _zz_DifftestDelayBundle_DifftestCsrRstat_2_2 <= _zz_DifftestDelayBundle_DifftestCsrRstat_2;
    _zz_DifftestDelayBundle_DifftestCsrRstat_3_2 <= _zz_DifftestDelayBundle_DifftestCsrRstat_3;
    _zz_DifftestDelayBundle_DifftestCsrRstat_4_2 <= _zz_DifftestDelayBundle_DifftestCsrRstat_4;
    _zz_DifftestDelayBundle_DifftestCsrData_0_2 <= _zz_DifftestDelayBundle_DifftestCsrData_0;
    _zz_DifftestDelayBundle_DifftestCsrData_1_2 <= _zz_DifftestDelayBundle_DifftestCsrData_1;
    _zz_DifftestDelayBundle_DifftestCsrData_2_2 <= _zz_DifftestDelayBundle_DifftestCsrData_2;
    _zz_DifftestDelayBundle_DifftestCsrData_3_2 <= _zz_DifftestDelayBundle_DifftestCsrData_3;
    _zz_DifftestDelayBundle_DifftestCsrData_4_2 <= _zz_DifftestDelayBundle_DifftestCsrData_4;
    _zz_DifftestDelayBundle_DifftestExcpEventExcpValid_2 <= _zz_DifftestDelayBundle_DifftestExcpEventExcpValid;
    _zz_DifftestDelayBundle_DifftestExcpEventEret_2 <= _zz_DifftestDelayBundle_DifftestExcpEventEret;
    _zz_DifftestDelayBundle_DifftestExcpEventIntrNO_2 <= _zz_DifftestDelayBundle_DifftestExcpEventIntrNO;
    _zz_DifftestDelayBundle_DifftestExcpEventCause_2 <= _zz_DifftestDelayBundle_DifftestExcpEventCause;
    _zz_DifftestDelayBundle_DifftestExcpEventEPC_2 <= _zz_DifftestDelayBundle_DifftestExcpEventEPC;
    _zz_DifftestDelayBundle_DifftestExcpEventInst_2 <= _zz_DifftestDelayBundle_DifftestExcpEventInst;
    _zz_DifftestDelayBundle_DifftestStoreEventValid_2 <= _zz_DifftestDelayBundle_DifftestStoreEventValid;
    _zz_DifftestDelayBundle_DifftestStoreEventPAddr_2 <= _zz_DifftestDelayBundle_DifftestStoreEventPAddr;
    _zz_DifftestDelayBundle_DifftestStoreEventVAddr_2 <= _zz_DifftestDelayBundle_DifftestStoreEventVAddr;
    _zz_DifftestDelayBundle_DifftestStoreEventData_2 <= _zz_DifftestDelayBundle_DifftestStoreEventData;
    _zz_DifftestDelayBundle_DifftestLoadEventValid_2 <= _zz_DifftestDelayBundle_DifftestLoadEventValid;
    _zz_DifftestDelayBundle_DifftestLoadEventPAddr_2 <= _zz_DifftestDelayBundle_DifftestLoadEventPAddr;
    _zz_DifftestDelayBundle_DifftestLoadEventVAddr_2 <= _zz_DifftestDelayBundle_DifftestLoadEventVAddr;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_0_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitIndex_0_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_1_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitIndex_1_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_2_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitIndex_2_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_3_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitIndex_3_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitIndex_4_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitIndex_4_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_0_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitValid_0_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_1_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitValid_1_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_2_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitValid_2_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_3_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitValid_3_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitValid_4_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitValid_4_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_0_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitPC_0_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_1_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitPC_1_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_2_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitPC_2_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_3_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitPC_3_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitPC_4_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitPC_4_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_0_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitInstr_0_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_1_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitInstr_1_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_2_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitInstr_2_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_3_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitInstr_3_2;
    _zz_DifftestDelayBundle_DifftestInstrCommitInstr_4_1 <= _zz_DifftestDelayBundle_DifftestInstrCommitInstr_4_2;
    _zz_DifftestDelayBundle_DifftestSkip_0_1 <= _zz_DifftestDelayBundle_DifftestSkip_0_2;
    _zz_DifftestDelayBundle_DifftestSkip_1_1 <= _zz_DifftestDelayBundle_DifftestSkip_1_2;
    _zz_DifftestDelayBundle_DifftestSkip_2_1 <= _zz_DifftestDelayBundle_DifftestSkip_2_2;
    _zz_DifftestDelayBundle_DifftestSkip_3_1 <= _zz_DifftestDelayBundle_DifftestSkip_3_2;
    _zz_DifftestDelayBundle_DifftestSkip_4_1 <= _zz_DifftestDelayBundle_DifftestSkip_4_2;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_0_1 <= _zz_DifftestDelayBundle_DifftestIsTlbFill_0_2;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_1_1 <= _zz_DifftestDelayBundle_DifftestIsTlbFill_1_2;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_2_1 <= _zz_DifftestDelayBundle_DifftestIsTlbFill_2_2;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_3_1 <= _zz_DifftestDelayBundle_DifftestIsTlbFill_3_2;
    _zz_DifftestDelayBundle_DifftestIsTlbFill_4_1 <= _zz_DifftestDelayBundle_DifftestIsTlbFill_4_2;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_0_1 <= _zz_DifftestDelayBundle_DifftestTlbFillIndex_0_2;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_1_1 <= _zz_DifftestDelayBundle_DifftestTlbFillIndex_1_2;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_2_1 <= _zz_DifftestDelayBundle_DifftestTlbFillIndex_2_2;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_3_1 <= _zz_DifftestDelayBundle_DifftestTlbFillIndex_3_2;
    _zz_DifftestDelayBundle_DifftestTlbFillIndex_4_1 <= _zz_DifftestDelayBundle_DifftestTlbFillIndex_4_2;
    _zz_DifftestDelayBundle_DifftestIsCount_0_1 <= _zz_DifftestDelayBundle_DifftestIsCount_0_2;
    _zz_DifftestDelayBundle_DifftestIsCount_1_1 <= _zz_DifftestDelayBundle_DifftestIsCount_1_2;
    _zz_DifftestDelayBundle_DifftestIsCount_2_1 <= _zz_DifftestDelayBundle_DifftestIsCount_2_2;
    _zz_DifftestDelayBundle_DifftestIsCount_3_1 <= _zz_DifftestDelayBundle_DifftestIsCount_3_2;
    _zz_DifftestDelayBundle_DifftestIsCount_4_1 <= _zz_DifftestDelayBundle_DifftestIsCount_4_2;
    _zz_DifftestDelayBundle_DifftestCount_0_1 <= _zz_DifftestDelayBundle_DifftestCount_0_2;
    _zz_DifftestDelayBundle_DifftestCount_1_1 <= _zz_DifftestDelayBundle_DifftestCount_1_2;
    _zz_DifftestDelayBundle_DifftestCount_2_1 <= _zz_DifftestDelayBundle_DifftestCount_2_2;
    _zz_DifftestDelayBundle_DifftestCount_3_1 <= _zz_DifftestDelayBundle_DifftestCount_3_2;
    _zz_DifftestDelayBundle_DifftestCount_4_1 <= _zz_DifftestDelayBundle_DifftestCount_4_2;
    _zz_DifftestDelayBundle_DifftestWen_0_1 <= _zz_DifftestDelayBundle_DifftestWen_0_2;
    _zz_DifftestDelayBundle_DifftestWen_1_1 <= _zz_DifftestDelayBundle_DifftestWen_1_2;
    _zz_DifftestDelayBundle_DifftestWen_2_1 <= _zz_DifftestDelayBundle_DifftestWen_2_2;
    _zz_DifftestDelayBundle_DifftestWen_3_1 <= _zz_DifftestDelayBundle_DifftestWen_3_2;
    _zz_DifftestDelayBundle_DifftestWen_4_1 <= _zz_DifftestDelayBundle_DifftestWen_4_2;
    _zz_DifftestDelayBundle_DifftestWdest_0_1 <= _zz_DifftestDelayBundle_DifftestWdest_0_2;
    _zz_DifftestDelayBundle_DifftestWdest_1_1 <= _zz_DifftestDelayBundle_DifftestWdest_1_2;
    _zz_DifftestDelayBundle_DifftestWdest_2_1 <= _zz_DifftestDelayBundle_DifftestWdest_2_2;
    _zz_DifftestDelayBundle_DifftestWdest_3_1 <= _zz_DifftestDelayBundle_DifftestWdest_3_2;
    _zz_DifftestDelayBundle_DifftestWdest_4_1 <= _zz_DifftestDelayBundle_DifftestWdest_4_2;
    _zz_DifftestDelayBundle_DifftestWdata_0_1 <= _zz_DifftestDelayBundle_DifftestWdata_0_2;
    _zz_DifftestDelayBundle_DifftestWdata_1_1 <= _zz_DifftestDelayBundle_DifftestWdata_1_2;
    _zz_DifftestDelayBundle_DifftestWdata_2_1 <= _zz_DifftestDelayBundle_DifftestWdata_2_2;
    _zz_DifftestDelayBundle_DifftestWdata_3_1 <= _zz_DifftestDelayBundle_DifftestWdata_3_2;
    _zz_DifftestDelayBundle_DifftestWdata_4_1 <= _zz_DifftestDelayBundle_DifftestWdata_4_2;
    _zz_DifftestDelayBundle_DifftestCsrRstat_0_1 <= _zz_DifftestDelayBundle_DifftestCsrRstat_0_2;
    _zz_DifftestDelayBundle_DifftestCsrRstat_1_1 <= _zz_DifftestDelayBundle_DifftestCsrRstat_1_2;
    _zz_DifftestDelayBundle_DifftestCsrRstat_2_1 <= _zz_DifftestDelayBundle_DifftestCsrRstat_2_2;
    _zz_DifftestDelayBundle_DifftestCsrRstat_3_1 <= _zz_DifftestDelayBundle_DifftestCsrRstat_3_2;
    _zz_DifftestDelayBundle_DifftestCsrRstat_4_1 <= _zz_DifftestDelayBundle_DifftestCsrRstat_4_2;
    _zz_DifftestDelayBundle_DifftestCsrData_0_1 <= _zz_DifftestDelayBundle_DifftestCsrData_0_2;
    _zz_DifftestDelayBundle_DifftestCsrData_1_1 <= _zz_DifftestDelayBundle_DifftestCsrData_1_2;
    _zz_DifftestDelayBundle_DifftestCsrData_2_1 <= _zz_DifftestDelayBundle_DifftestCsrData_2_2;
    _zz_DifftestDelayBundle_DifftestCsrData_3_1 <= _zz_DifftestDelayBundle_DifftestCsrData_3_2;
    _zz_DifftestDelayBundle_DifftestCsrData_4_1 <= _zz_DifftestDelayBundle_DifftestCsrData_4_2;
    _zz_DifftestDelayBundle_DifftestExcpEventExcpValid_1 <= _zz_DifftestDelayBundle_DifftestExcpEventExcpValid_2;
    _zz_DifftestDelayBundle_DifftestExcpEventEret_1 <= _zz_DifftestDelayBundle_DifftestExcpEventEret_2;
    _zz_DifftestDelayBundle_DifftestExcpEventIntrNO_1 <= _zz_DifftestDelayBundle_DifftestExcpEventIntrNO_2;
    _zz_DifftestDelayBundle_DifftestExcpEventCause_1 <= _zz_DifftestDelayBundle_DifftestExcpEventCause_2;
    _zz_DifftestDelayBundle_DifftestExcpEventEPC_1 <= _zz_DifftestDelayBundle_DifftestExcpEventEPC_2;
    _zz_DifftestDelayBundle_DifftestExcpEventInst_1 <= _zz_DifftestDelayBundle_DifftestExcpEventInst_2;
    _zz_DifftestDelayBundle_DifftestStoreEventValid_1 <= _zz_DifftestDelayBundle_DifftestStoreEventValid_2;
    _zz_DifftestDelayBundle_DifftestStoreEventPAddr_1 <= _zz_DifftestDelayBundle_DifftestStoreEventPAddr_2;
    _zz_DifftestDelayBundle_DifftestStoreEventVAddr_1 <= _zz_DifftestDelayBundle_DifftestStoreEventVAddr_2;
    _zz_DifftestDelayBundle_DifftestStoreEventData_1 <= _zz_DifftestDelayBundle_DifftestStoreEventData_2;
    _zz_DifftestDelayBundle_DifftestLoadEventValid_1 <= _zz_DifftestDelayBundle_DifftestLoadEventValid_2;
    _zz_DifftestDelayBundle_DifftestLoadEventPAddr_1 <= _zz_DifftestDelayBundle_DifftestLoadEventPAddr_2;
    _zz_DifftestDelayBundle_DifftestLoadEventVAddr_1 <= _zz_DifftestDelayBundle_DifftestLoadEventVAddr_2;
  end


endmodule

//CommitLogic_4 replaced by CommitLogic

//CommitLogic_3 replaced by CommitLogic

//CommitLogic_2 replaced by CommitLogic

//CommitLogic_1 replaced by CommitLogic

module CommitLogic (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [4:0]    io_input_payload_robIdx,
  input  wire [31:0]   io_input_payload_data,
  input  wire [5:0]    io_input_payload_prd,
  input  wire [31:0]   io_input_payload_branchResult_targetPC,
  input  wire          io_input_payload_branchResult_branchResult,
  input  wire          io_input_payload_branchResult_predictFail,
  input  wire          io_input_payload_exceptionInfo_exception,
  input  wire [5:0]    io_input_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_input_payload_exceptionInfo_eSubCode,
  output wire [5:0]    io_srat_prd,
  output wire          io_srat_wen,
  output wire [4:0]    io_rob_robIdx,
  output wire [31:0]   io_rob_branchResult_targetPC,
  output wire          io_rob_branchResult_branchResult,
  output wire          io_rob_branchResult_predictFail,
  output wire          io_rob_exceptionInfo_exception,
  output wire [5:0]    io_rob_exceptionInfo_eCode,
  output wire [0:0]    io_rob_exceptionInfo_eSubCode,
  output wire          io_rob_valid,
  output wire [5:0]    io_prf_idx,
  output wire [31:0]   io_prf_data,
  output wire          io_forward_valid,
  output wire [5:0]    io_forward_payload_idx,
  output wire [31:0]   io_forward_payload_payload
);


  assign io_input_ready = 1'b1;
  assign io_srat_prd = io_input_payload_prd;
  assign io_srat_wen = io_input_valid;
  assign io_rob_robIdx = io_input_payload_robIdx;
  assign io_rob_branchResult_targetPC = io_input_payload_branchResult_targetPC;
  assign io_rob_branchResult_branchResult = io_input_payload_branchResult_branchResult;
  assign io_rob_branchResult_predictFail = io_input_payload_branchResult_predictFail;
  assign io_rob_exceptionInfo_exception = io_input_payload_exceptionInfo_exception;
  assign io_rob_exceptionInfo_eCode = io_input_payload_exceptionInfo_eCode;
  assign io_rob_exceptionInfo_eSubCode = io_input_payload_exceptionInfo_eSubCode;
  assign io_rob_valid = io_input_valid;
  assign io_prf_idx = (io_input_valid ? io_input_payload_prd : 6'h00);
  assign io_prf_data = io_input_payload_data;
  assign io_forward_valid = (io_input_valid && (io_input_payload_prd != 6'h00));
  assign io_forward_payload_idx = io_input_payload_prd;
  assign io_forward_payload_payload = io_input_payload_data;

endmodule

module DIVU (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [31:0]   io_input_payload_src1,
  input  wire [31:0]   io_input_payload_src2,
  input  wire [4:0]    io_input_payload_robIdx,
  input  wire [31:0]   io_input_payload_branchResult_targetPC,
  input  wire          io_input_payload_branchResult_branchResult,
  input  wire          io_input_payload_branchResult_predictFail,
  input  wire          io_input_payload_exceptionInfo_exception,
  input  wire [5:0]    io_input_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_input_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_payload_pc,
  input  wire [5:0]    io_input_payload_prd,
  input  wire [1:0]    io_input_payload_uop_divuOp,
  output reg           io_output_valid,
  input  wire          io_output_ready,
  output wire [4:0]    io_output_payload_robIdx,
  output reg  [31:0]   io_output_payload_data,
  output wire [5:0]    io_output_payload_prd,
  output wire [31:0]   io_output_payload_branchResult_targetPC,
  output wire          io_output_payload_branchResult_branchResult,
  output wire          io_output_payload_branchResult_predictFail,
  output wire          io_output_payload_exceptionInfo_exception,
  output wire [5:0]    io_output_payload_exceptionInfo_eCode,
  output wire [0:0]    io_output_payload_exceptionInfo_eSubCode,
  input  wire          aclk,
  input  wire          cpuClockingArea_areaFlushReset_newReset
);
  localparam DIVUOp_div = 2'd0;
  localparam DIVUOp_divu = 2'd1;
  localparam DIVUOp_mod_1 = 2'd2;
  localparam DIVUOp_modu = 2'd3;

  wire       [5:0]    _zz_counter_valueNext;
  wire       [0:0]    _zz_counter_valueNext_1;
  wire       [31:0]   _zz_io_output_payload_data;
  wire       [31:0]   _zz_io_output_payload_data_1;
  wire       [31:0]   _zz_io_output_payload_data_2;
  wire       [31:0]   _zz_io_output_payload_data_3;
  wire       [31:0]   _zz_io_output_payload_data_4;
  wire       [31:0]   _zz_io_output_payload_data_5;
  reg                 block_1;
  reg                 counter_willIncrement;
  wire                counter_willClear;
  reg        [5:0]    counter_valueNext;
  reg        [5:0]    counter_value;
  wire                counter_willOverflowIfInc;
  wire                counter_willOverflow;
  wire                io_input_fire;
  wire                when_DIVU_l26;
  `ifndef SYNTHESIS
  reg [39:0] io_input_payload_uop_divuOp_string;
  `endif


  assign _zz_counter_valueNext_1 = counter_willIncrement;
  assign _zz_counter_valueNext = {5'd0, _zz_counter_valueNext_1};
  assign _zz_io_output_payload_data = ($signed(_zz_io_output_payload_data_1) / $signed(_zz_io_output_payload_data_2));
  assign _zz_io_output_payload_data_1 = io_input_payload_src1;
  assign _zz_io_output_payload_data_2 = io_input_payload_src2;
  assign _zz_io_output_payload_data_3 = ($signed(_zz_io_output_payload_data_4) % $signed(_zz_io_output_payload_data_5));
  assign _zz_io_output_payload_data_4 = io_input_payload_src1;
  assign _zz_io_output_payload_data_5 = io_input_payload_src2;
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_uop_divuOp)
      DIVUOp_div : io_input_payload_uop_divuOp_string = "div  ";
      DIVUOp_divu : io_input_payload_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : io_input_payload_uop_divuOp_string = "mod_1";
      DIVUOp_modu : io_input_payload_uop_divuOp_string = "modu ";
      default : io_input_payload_uop_divuOp_string = "?????";
    endcase
  end
  `endif

  always @(*) begin
    counter_willIncrement = 1'b0;
    if(block_1) begin
      counter_willIncrement = 1'b1;
    end
  end

  assign counter_willClear = 1'b0;
  assign counter_willOverflowIfInc = (counter_value == 6'h20);
  assign counter_willOverflow = (counter_willOverflowIfInc && counter_willIncrement);
  always @(*) begin
    if(counter_willOverflow) begin
      counter_valueNext = 6'h00;
    end else begin
      counter_valueNext = (counter_value + _zz_counter_valueNext);
    end
    if(counter_willClear) begin
      counter_valueNext = 6'h00;
    end
  end

  assign io_input_ready = (! block_1);
  always @(*) begin
    io_output_valid = 1'b0;
    if(when_DIVU_l26) begin
      io_output_valid = 1'b1;
    end
  end

  assign io_input_fire = (io_input_valid && io_input_ready);
  assign when_DIVU_l26 = (counter_willOverflowIfInc || (block_1 && io_input_payload_exceptionInfo_exception));
  assign io_output_payload_robIdx = io_input_payload_robIdx;
  assign io_output_payload_prd = io_input_payload_prd;
  assign io_output_payload_branchResult_targetPC = io_input_payload_branchResult_targetPC;
  assign io_output_payload_branchResult_branchResult = io_input_payload_branchResult_branchResult;
  assign io_output_payload_branchResult_predictFail = io_input_payload_branchResult_predictFail;
  assign io_output_payload_exceptionInfo_exception = io_input_payload_exceptionInfo_exception;
  assign io_output_payload_exceptionInfo_eCode = io_input_payload_exceptionInfo_eCode;
  assign io_output_payload_exceptionInfo_eSubCode = io_input_payload_exceptionInfo_eSubCode;
  always @(*) begin
    case(io_input_payload_uop_divuOp)
      DIVUOp_div : begin
        io_output_payload_data = _zz_io_output_payload_data;
      end
      DIVUOp_divu : begin
        io_output_payload_data = (io_input_payload_src1 / io_input_payload_src2);
      end
      DIVUOp_mod_1 : begin
        io_output_payload_data = _zz_io_output_payload_data_3;
      end
      default : begin
        io_output_payload_data = (io_input_payload_src1 % io_input_payload_src2);
      end
    endcase
  end

  always @(posedge aclk) begin
    if(!cpuClockingArea_areaFlushReset_newReset) begin
      block_1 <= 1'b0;
      counter_value <= 6'h00;
    end else begin
      counter_value <= counter_valueNext;
      block_1 <= block_1;
      if(io_input_fire) begin
        block_1 <= 1'b1;
      end
      if(when_DIVU_l26) begin
        block_1 <= 1'b0;
      end
    end
  end


endmodule

module MULU (
  input  wire          io_input_valid,
  output reg           io_input_ready,
  input  wire [31:0]   io_input_payload_src1,
  input  wire [31:0]   io_input_payload_src2,
  input  wire [4:0]    io_input_payload_robIdx,
  input  wire [31:0]   io_input_payload_branchResult_targetPC,
  input  wire          io_input_payload_branchResult_branchResult,
  input  wire          io_input_payload_branchResult_predictFail,
  input  wire          io_input_payload_exceptionInfo_exception,
  input  wire [5:0]    io_input_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_input_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_payload_pc,
  input  wire [5:0]    io_input_payload_prd,
  input  wire [1:0]    io_input_payload_uop_muluOp,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [4:0]    io_output_payload_robIdx,
  output wire [31:0]   io_output_payload_data,
  output wire [5:0]    io_output_payload_prd,
  output wire [31:0]   io_output_payload_branchResult_targetPC,
  output wire          io_output_payload_branchResult_branchResult,
  output wire          io_output_payload_branchResult_predictFail,
  output wire          io_output_payload_exceptionInfo_exception,
  output wire [5:0]    io_output_payload_exceptionInfo_eCode,
  output wire [0:0]    io_output_payload_exceptionInfo_eSubCode,
  output wire          io_forward_valid,
  output wire [5:0]    io_forward_payload_idx,
  output wire [31:0]   io_forward_payload_payload,
  output wire          io_wakeOut_0_valid,
  output wire [5:0]    io_wakeOut_0_payload,
  output wire          io_wakeOut_1_valid,
  output wire [5:0]    io_wakeOut_1_payload,
  output wire          io_wakeOut_2_valid,
  output wire [5:0]    io_wakeOut_2_payload,
  input  wire          aclk,
  input  wire          cpuClockingArea_areaFlushReset_newReset
);
  localparam MULUOp_mullo = 2'd0;
  localparam MULUOp_mulhi = 2'd1;
  localparam MULUOp_mulhiu = 2'd2;

  wire       [31:0]   _zz_ress;
  wire       [31:0]   _zz_ress_1;
  wire       [31:0]   _zz_res;
  wire                stage12_valid;
  reg                 stage12_ready;
  wire       [31:0]   stage12_payload_src1;
  wire       [31:0]   stage12_payload_src2;
  wire       [4:0]    stage12_payload_robIdx;
  wire       [31:0]   stage12_payload_branchResult_targetPC;
  wire                stage12_payload_branchResult_branchResult;
  wire                stage12_payload_branchResult_predictFail;
  wire                stage12_payload_exceptionInfo_exception;
  wire       [5:0]    stage12_payload_exceptionInfo_eCode;
  wire       [0:0]    stage12_payload_exceptionInfo_eSubCode;
  wire       [31:0]   stage12_payload_pc;
  wire       [5:0]    stage12_payload_prd;
  wire       [1:0]    stage12_payload_uop_muluOp;
  wire                io_input_m2sPipe_valid;
  wire                io_input_m2sPipe_ready;
  wire       [31:0]   io_input_m2sPipe_payload_src1;
  wire       [31:0]   io_input_m2sPipe_payload_src2;
  wire       [4:0]    io_input_m2sPipe_payload_robIdx;
  wire       [31:0]   io_input_m2sPipe_payload_branchResult_targetPC;
  wire                io_input_m2sPipe_payload_branchResult_branchResult;
  wire                io_input_m2sPipe_payload_branchResult_predictFail;
  wire                io_input_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    io_input_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    io_input_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   io_input_m2sPipe_payload_pc;
  wire       [5:0]    io_input_m2sPipe_payload_prd;
  wire       [1:0]    io_input_m2sPipe_payload_uop_muluOp;
  reg                 io_input_rValid;
  reg        [31:0]   io_input_rData_src1;
  reg        [31:0]   io_input_rData_src2;
  reg        [4:0]    io_input_rData_robIdx;
  reg        [31:0]   io_input_rData_branchResult_targetPC;
  reg                 io_input_rData_branchResult_branchResult;
  reg                 io_input_rData_branchResult_predictFail;
  reg                 io_input_rData_exceptionInfo_exception;
  reg        [5:0]    io_input_rData_exceptionInfo_eCode;
  reg        [0:0]    io_input_rData_exceptionInfo_eSubCode;
  reg        [31:0]   io_input_rData_pc;
  reg        [5:0]    io_input_rData_prd;
  reg        [1:0]    io_input_rData_uop_muluOp;
  wire                when_Stream_l369;
  wire                stage23_valid;
  wire                stage23_ready;
  wire       [31:0]   stage23_payload_src1;
  wire       [31:0]   stage23_payload_src2;
  wire       [4:0]    stage23_payload_robIdx;
  wire       [31:0]   stage23_payload_branchResult_targetPC;
  wire                stage23_payload_branchResult_branchResult;
  wire                stage23_payload_branchResult_predictFail;
  wire                stage23_payload_exceptionInfo_exception;
  wire       [5:0]    stage23_payload_exceptionInfo_eCode;
  wire       [0:0]    stage23_payload_exceptionInfo_eSubCode;
  wire       [31:0]   stage23_payload_pc;
  wire       [5:0]    stage23_payload_prd;
  wire       [1:0]    stage23_payload_uop_muluOp;
  wire                stage12_m2sPipe_valid;
  wire                stage12_m2sPipe_ready;
  wire       [31:0]   stage12_m2sPipe_payload_src1;
  wire       [31:0]   stage12_m2sPipe_payload_src2;
  wire       [4:0]    stage12_m2sPipe_payload_robIdx;
  wire       [31:0]   stage12_m2sPipe_payload_branchResult_targetPC;
  wire                stage12_m2sPipe_payload_branchResult_branchResult;
  wire                stage12_m2sPipe_payload_branchResult_predictFail;
  wire                stage12_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    stage12_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    stage12_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   stage12_m2sPipe_payload_pc;
  wire       [5:0]    stage12_m2sPipe_payload_prd;
  wire       [1:0]    stage12_m2sPipe_payload_uop_muluOp;
  reg                 stage12_rValid;
  reg        [31:0]   stage12_rData_src1;
  reg        [31:0]   stage12_rData_src2;
  reg        [4:0]    stage12_rData_robIdx;
  reg        [31:0]   stage12_rData_branchResult_targetPC;
  reg                 stage12_rData_branchResult_branchResult;
  reg                 stage12_rData_branchResult_predictFail;
  reg                 stage12_rData_exceptionInfo_exception;
  reg        [5:0]    stage12_rData_exceptionInfo_eCode;
  reg        [0:0]    stage12_rData_exceptionInfo_eSubCode;
  reg        [31:0]   stage12_rData_pc;
  reg        [5:0]    stage12_rData_prd;
  reg        [1:0]    stage12_rData_uop_muluOp;
  wire                when_Stream_l369_1;
  wire       [63:0]   resu;
  wire       [63:0]   ress;
  reg        [31:0]   res;
  `ifndef SYNTHESIS
  reg [47:0] io_input_payload_uop_muluOp_string;
  reg [47:0] stage12_payload_uop_muluOp_string;
  reg [47:0] io_input_m2sPipe_payload_uop_muluOp_string;
  reg [47:0] io_input_rData_uop_muluOp_string;
  reg [47:0] stage23_payload_uop_muluOp_string;
  reg [47:0] stage12_m2sPipe_payload_uop_muluOp_string;
  reg [47:0] stage12_rData_uop_muluOp_string;
  `endif


  assign _zz_ress = stage23_payload_src1;
  assign _zz_ress_1 = stage23_payload_src2;
  assign _zz_res = ress[63 : 32];
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_uop_muluOp)
      MULUOp_mullo : io_input_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : io_input_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : io_input_payload_uop_muluOp_string = "mulhiu";
      default : io_input_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(stage12_payload_uop_muluOp)
      MULUOp_mullo : stage12_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : stage12_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : stage12_payload_uop_muluOp_string = "mulhiu";
      default : stage12_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_input_m2sPipe_payload_uop_muluOp)
      MULUOp_mullo : io_input_m2sPipe_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : io_input_m2sPipe_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : io_input_m2sPipe_payload_uop_muluOp_string = "mulhiu";
      default : io_input_m2sPipe_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_input_rData_uop_muluOp)
      MULUOp_mullo : io_input_rData_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : io_input_rData_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : io_input_rData_uop_muluOp_string = "mulhiu";
      default : io_input_rData_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(stage23_payload_uop_muluOp)
      MULUOp_mullo : stage23_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : stage23_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : stage23_payload_uop_muluOp_string = "mulhiu";
      default : stage23_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(stage12_m2sPipe_payload_uop_muluOp)
      MULUOp_mullo : stage12_m2sPipe_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : stage12_m2sPipe_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : stage12_m2sPipe_payload_uop_muluOp_string = "mulhiu";
      default : stage12_m2sPipe_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(stage12_rData_uop_muluOp)
      MULUOp_mullo : stage12_rData_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : stage12_rData_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : stage12_rData_uop_muluOp_string = "mulhiu";
      default : stage12_rData_uop_muluOp_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    io_input_ready = io_input_m2sPipe_ready;
    if(when_Stream_l369) begin
      io_input_ready = 1'b1;
    end
  end

  assign when_Stream_l369 = (! io_input_m2sPipe_valid);
  assign io_input_m2sPipe_valid = io_input_rValid;
  assign io_input_m2sPipe_payload_src1 = io_input_rData_src1;
  assign io_input_m2sPipe_payload_src2 = io_input_rData_src2;
  assign io_input_m2sPipe_payload_robIdx = io_input_rData_robIdx;
  assign io_input_m2sPipe_payload_branchResult_targetPC = io_input_rData_branchResult_targetPC;
  assign io_input_m2sPipe_payload_branchResult_branchResult = io_input_rData_branchResult_branchResult;
  assign io_input_m2sPipe_payload_branchResult_predictFail = io_input_rData_branchResult_predictFail;
  assign io_input_m2sPipe_payload_exceptionInfo_exception = io_input_rData_exceptionInfo_exception;
  assign io_input_m2sPipe_payload_exceptionInfo_eCode = io_input_rData_exceptionInfo_eCode;
  assign io_input_m2sPipe_payload_exceptionInfo_eSubCode = io_input_rData_exceptionInfo_eSubCode;
  assign io_input_m2sPipe_payload_pc = io_input_rData_pc;
  assign io_input_m2sPipe_payload_prd = io_input_rData_prd;
  assign io_input_m2sPipe_payload_uop_muluOp = io_input_rData_uop_muluOp;
  assign stage12_valid = io_input_m2sPipe_valid;
  assign io_input_m2sPipe_ready = stage12_ready;
  assign stage12_payload_src1 = io_input_m2sPipe_payload_src1;
  assign stage12_payload_src2 = io_input_m2sPipe_payload_src2;
  assign stage12_payload_robIdx = io_input_m2sPipe_payload_robIdx;
  assign stage12_payload_branchResult_targetPC = io_input_m2sPipe_payload_branchResult_targetPC;
  assign stage12_payload_branchResult_branchResult = io_input_m2sPipe_payload_branchResult_branchResult;
  assign stage12_payload_branchResult_predictFail = io_input_m2sPipe_payload_branchResult_predictFail;
  assign stage12_payload_exceptionInfo_exception = io_input_m2sPipe_payload_exceptionInfo_exception;
  assign stage12_payload_exceptionInfo_eCode = io_input_m2sPipe_payload_exceptionInfo_eCode;
  assign stage12_payload_exceptionInfo_eSubCode = io_input_m2sPipe_payload_exceptionInfo_eSubCode;
  assign stage12_payload_pc = io_input_m2sPipe_payload_pc;
  assign stage12_payload_prd = io_input_m2sPipe_payload_prd;
  assign stage12_payload_uop_muluOp = io_input_m2sPipe_payload_uop_muluOp;
  always @(*) begin
    stage12_ready = stage12_m2sPipe_ready;
    if(when_Stream_l369_1) begin
      stage12_ready = 1'b1;
    end
  end

  assign when_Stream_l369_1 = (! stage12_m2sPipe_valid);
  assign stage12_m2sPipe_valid = stage12_rValid;
  assign stage12_m2sPipe_payload_src1 = stage12_rData_src1;
  assign stage12_m2sPipe_payload_src2 = stage12_rData_src2;
  assign stage12_m2sPipe_payload_robIdx = stage12_rData_robIdx;
  assign stage12_m2sPipe_payload_branchResult_targetPC = stage12_rData_branchResult_targetPC;
  assign stage12_m2sPipe_payload_branchResult_branchResult = stage12_rData_branchResult_branchResult;
  assign stage12_m2sPipe_payload_branchResult_predictFail = stage12_rData_branchResult_predictFail;
  assign stage12_m2sPipe_payload_exceptionInfo_exception = stage12_rData_exceptionInfo_exception;
  assign stage12_m2sPipe_payload_exceptionInfo_eCode = stage12_rData_exceptionInfo_eCode;
  assign stage12_m2sPipe_payload_exceptionInfo_eSubCode = stage12_rData_exceptionInfo_eSubCode;
  assign stage12_m2sPipe_payload_pc = stage12_rData_pc;
  assign stage12_m2sPipe_payload_prd = stage12_rData_prd;
  assign stage12_m2sPipe_payload_uop_muluOp = stage12_rData_uop_muluOp;
  assign stage23_valid = stage12_m2sPipe_valid;
  assign stage12_m2sPipe_ready = stage23_ready;
  assign stage23_payload_src1 = stage12_m2sPipe_payload_src1;
  assign stage23_payload_src2 = stage12_m2sPipe_payload_src2;
  assign stage23_payload_robIdx = stage12_m2sPipe_payload_robIdx;
  assign stage23_payload_branchResult_targetPC = stage12_m2sPipe_payload_branchResult_targetPC;
  assign stage23_payload_branchResult_branchResult = stage12_m2sPipe_payload_branchResult_branchResult;
  assign stage23_payload_branchResult_predictFail = stage12_m2sPipe_payload_branchResult_predictFail;
  assign stage23_payload_exceptionInfo_exception = stage12_m2sPipe_payload_exceptionInfo_exception;
  assign stage23_payload_exceptionInfo_eCode = stage12_m2sPipe_payload_exceptionInfo_eCode;
  assign stage23_payload_exceptionInfo_eSubCode = stage12_m2sPipe_payload_exceptionInfo_eSubCode;
  assign stage23_payload_pc = stage12_m2sPipe_payload_pc;
  assign stage23_payload_prd = stage12_m2sPipe_payload_prd;
  assign stage23_payload_uop_muluOp = stage12_m2sPipe_payload_uop_muluOp;
  assign resu = (stage23_payload_src1 * stage23_payload_src2);
  assign ress = ($signed(_zz_ress) * $signed(_zz_ress_1));
  assign io_forward_valid = (stage23_valid && (stage23_payload_prd != 6'h00));
  assign io_forward_payload_idx = stage23_payload_prd;
  assign io_forward_payload_payload = res;
  assign io_output_valid = stage23_valid;
  assign stage23_ready = io_output_ready;
  assign io_output_payload_robIdx = stage23_payload_robIdx;
  assign io_output_payload_data = res;
  assign io_output_payload_prd = stage23_payload_prd;
  assign io_output_payload_branchResult_targetPC = stage23_payload_branchResult_targetPC;
  assign io_output_payload_branchResult_branchResult = stage23_payload_branchResult_branchResult;
  assign io_output_payload_branchResult_predictFail = stage23_payload_branchResult_predictFail;
  assign io_output_payload_exceptionInfo_exception = stage23_payload_exceptionInfo_exception;
  assign io_output_payload_exceptionInfo_eCode = stage23_payload_exceptionInfo_eCode;
  assign io_output_payload_exceptionInfo_eSubCode = stage23_payload_exceptionInfo_eSubCode;
  always @(*) begin
    case(stage23_payload_uop_muluOp)
      MULUOp_mullo : begin
        res = resu[31 : 0];
      end
      MULUOp_mulhi : begin
        res = _zz_res;
      end
      default : begin
        res = resu[63 : 32];
      end
    endcase
  end

  assign io_wakeOut_0_valid = io_input_valid;
  assign io_wakeOut_0_payload = io_input_payload_prd;
  assign io_wakeOut_1_valid = stage12_valid;
  assign io_wakeOut_1_payload = stage12_payload_prd;
  assign io_wakeOut_2_valid = stage23_valid;
  assign io_wakeOut_2_payload = stage23_payload_prd;
  always @(posedge aclk) begin
    if(!cpuClockingArea_areaFlushReset_newReset) begin
      io_input_rValid <= 1'b0;
      stage12_rValid <= 1'b0;
    end else begin
      if(io_input_ready) begin
        io_input_rValid <= io_input_valid;
      end
      if(stage12_ready) begin
        stage12_rValid <= stage12_valid;
      end
    end
  end

  always @(posedge aclk) begin
    if(io_input_ready) begin
      io_input_rData_src1 <= io_input_payload_src1;
      io_input_rData_src2 <= io_input_payload_src2;
      io_input_rData_robIdx <= io_input_payload_robIdx;
      io_input_rData_branchResult_targetPC <= io_input_payload_branchResult_targetPC;
      io_input_rData_branchResult_branchResult <= io_input_payload_branchResult_branchResult;
      io_input_rData_branchResult_predictFail <= io_input_payload_branchResult_predictFail;
      io_input_rData_exceptionInfo_exception <= io_input_payload_exceptionInfo_exception;
      io_input_rData_exceptionInfo_eCode <= io_input_payload_exceptionInfo_eCode;
      io_input_rData_exceptionInfo_eSubCode <= io_input_payload_exceptionInfo_eSubCode;
      io_input_rData_pc <= io_input_payload_pc;
      io_input_rData_prd <= io_input_payload_prd;
      io_input_rData_uop_muluOp <= io_input_payload_uop_muluOp;
    end
    if(stage12_ready) begin
      stage12_rData_src1 <= stage12_payload_src1;
      stage12_rData_src2 <= stage12_payload_src2;
      stage12_rData_robIdx <= stage12_payload_robIdx;
      stage12_rData_branchResult_targetPC <= stage12_payload_branchResult_targetPC;
      stage12_rData_branchResult_branchResult <= stage12_payload_branchResult_branchResult;
      stage12_rData_branchResult_predictFail <= stage12_payload_branchResult_predictFail;
      stage12_rData_exceptionInfo_exception <= stage12_payload_exceptionInfo_exception;
      stage12_rData_exceptionInfo_eCode <= stage12_payload_exceptionInfo_eCode;
      stage12_rData_exceptionInfo_eSubCode <= stage12_payload_exceptionInfo_eSubCode;
      stage12_rData_pc <= stage12_payload_pc;
      stage12_rData_prd <= stage12_payload_prd;
      stage12_rData_uop_muluOp <= stage12_payload_uop_muluOp;
    end
  end


endmodule

module ALU_1 (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [31:0]   io_input_payload_src1,
  input  wire [31:0]   io_input_payload_src2,
  input  wire [31:0]   io_input_payload_src3,
  input  wire [31:0]   io_input_payload_src4,
  input  wire [4:0]    io_input_payload_robIdx,
  input  wire [31:0]   io_input_payload_branchInfo_predictPC,
  input  wire          io_input_payload_branchInfo_predictResult,
  input  wire          io_input_payload_exceptionInfo_exception,
  input  wire [5:0]    io_input_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_input_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_payload_pc,
  input  wire [5:0]    io_input_payload_prd,
  input  wire [3:0]    io_input_payload_uop_aluOp,
  input  wire [1:0]    io_input_payload_uop_bruOp,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [4:0]    io_output_payload_robIdx,
  output reg  [31:0]   io_output_payload_data,
  output wire [5:0]    io_output_payload_prd,
  output wire [31:0]   io_output_payload_branchResult_targetPC,
  output reg           io_output_payload_branchResult_branchResult,
  output wire          io_output_payload_branchResult_predictFail,
  output wire          io_output_payload_exceptionInfo_exception,
  output wire [5:0]    io_output_payload_exceptionInfo_eCode,
  output wire [0:0]    io_output_payload_exceptionInfo_eSubCode,
  output wire          io_forward_valid,
  output wire [5:0]    io_forward_payload_idx,
  output wire [31:0]   io_forward_payload_payload,
  output wire          io_wakeOut_valid,
  output wire [5:0]    io_wakeOut_payload
);
  localparam ALUOp_add = 4'd0;
  localparam ALUOp_sub = 4'd1;
  localparam ALUOp_slt = 4'd2;
  localparam ALUOp_sltu = 4'd3;
  localparam ALUOp_eq = 4'd4;
  localparam ALUOp_nor_1 = 4'd5;
  localparam ALUOp_and_1 = 4'd6;
  localparam ALUOp_or_1 = 4'd7;
  localparam ALUOp_xor_1 = 4'd8;
  localparam ALUOp_sll_1 = 4'd9;
  localparam ALUOp_srl_1 = 4'd10;
  localparam ALUOp_sra_1 = 4'd11;
  localparam ALUOp_passa = 4'd12;
  localparam ALUOp_passb = 4'd13;
  localparam BRUOp_nop = 2'd0;
  localparam BRUOp_add = 2'd1;
  localparam BRUOp_cadd = 2'd2;
  localparam BRUOp_ncadd = 2'd3;

  wire       [31:0]   _zz_slt;
  wire       [31:0]   _zz_slt_1;
  wire       [31:0]   _zz_sra_1;
  wire       [31:0]   _zz_sra_1_1;
  wire       [31:0]   add;
  wire       [31:0]   sub;
  wire       [0:0]    slt;
  wire       [0:0]    sltu;
  wire       [0:0]    eq;
  wire       [31:0]   nor_1;
  wire       [31:0]   and_1;
  wire       [31:0]   or_1;
  wire       [31:0]   xor_1;
  wire       [31:0]   sll_1;
  wire       [31:0]   srl_1;
  wire       [31:0]   sra_1;
  `ifndef SYNTHESIS
  reg [39:0] io_input_payload_uop_aluOp_string;
  reg [39:0] io_input_payload_uop_bruOp_string;
  `endif


  assign _zz_slt = io_input_payload_src1;
  assign _zz_slt_1 = io_input_payload_src2;
  assign _zz_sra_1 = ($signed(_zz_sra_1_1) >>> io_input_payload_src2[4 : 0]);
  assign _zz_sra_1_1 = io_input_payload_src1;
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_uop_aluOp)
      ALUOp_add : io_input_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_input_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_input_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_input_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_input_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_input_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_input_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_input_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_input_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_input_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_input_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_input_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_input_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_input_payload_uop_aluOp_string = "passb";
      default : io_input_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_input_payload_uop_bruOp)
      BRUOp_nop : io_input_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_input_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_input_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_input_payload_uop_bruOp_string = "ncadd";
      default : io_input_payload_uop_bruOp_string = "?????";
    endcase
  end
  `endif

  assign io_input_ready = io_output_ready;
  assign io_output_valid = io_input_valid;
  assign io_output_payload_robIdx = io_input_payload_robIdx;
  assign io_output_payload_prd = io_input_payload_prd;
  assign io_output_payload_exceptionInfo_exception = io_input_payload_exceptionInfo_exception;
  assign io_output_payload_exceptionInfo_eCode = io_input_payload_exceptionInfo_eCode;
  assign io_output_payload_exceptionInfo_eSubCode = io_input_payload_exceptionInfo_eSubCode;
  assign io_forward_valid = (io_input_valid && (io_input_payload_prd != 6'h00));
  assign io_forward_payload_idx = io_input_payload_prd;
  assign io_forward_payload_payload = io_output_payload_data;
  assign io_wakeOut_valid = io_input_valid;
  assign io_wakeOut_payload = io_input_payload_prd;
  assign add = (io_input_payload_src1 + io_input_payload_src2);
  assign sub = (io_input_payload_src1 - io_input_payload_src2);
  assign slt = ($signed(_zz_slt) < $signed(_zz_slt_1));
  assign sltu = (io_input_payload_src1 < io_input_payload_src2);
  assign eq = (io_input_payload_src1 == io_input_payload_src2);
  assign nor_1 = (~ (io_input_payload_src1 | io_input_payload_src2));
  assign and_1 = (io_input_payload_src1 & io_input_payload_src2);
  assign or_1 = (io_input_payload_src1 | io_input_payload_src2);
  assign xor_1 = (io_input_payload_src1 ^ io_input_payload_src2);
  assign sll_1 = (io_input_payload_src1 <<< io_input_payload_src2[4 : 0]);
  assign srl_1 = (io_input_payload_src1 >>> io_input_payload_src2[4 : 0]);
  assign sra_1 = _zz_sra_1;
  always @(*) begin
    case(io_input_payload_uop_aluOp)
      ALUOp_add : begin
        io_output_payload_data = add;
      end
      ALUOp_sub : begin
        io_output_payload_data = sub;
      end
      ALUOp_slt : begin
        io_output_payload_data = {31'd0, slt};
      end
      ALUOp_sltu : begin
        io_output_payload_data = {31'd0, sltu};
      end
      ALUOp_eq : begin
        io_output_payload_data = {31'd0, eq};
      end
      ALUOp_nor_1 : begin
        io_output_payload_data = nor_1;
      end
      ALUOp_and_1 : begin
        io_output_payload_data = and_1;
      end
      ALUOp_or_1 : begin
        io_output_payload_data = or_1;
      end
      ALUOp_xor_1 : begin
        io_output_payload_data = xor_1;
      end
      ALUOp_sll_1 : begin
        io_output_payload_data = sll_1;
      end
      ALUOp_srl_1 : begin
        io_output_payload_data = srl_1;
      end
      ALUOp_sra_1 : begin
        io_output_payload_data = sra_1;
      end
      ALUOp_passa : begin
        io_output_payload_data = io_input_payload_src1;
      end
      default : begin
        io_output_payload_data = io_input_payload_src2;
      end
    endcase
  end

  assign io_output_payload_branchResult_targetPC = (io_input_payload_src3 + io_input_payload_src4);
  assign io_output_payload_branchResult_predictFail = (((io_output_payload_branchResult_targetPC != io_input_payload_branchInfo_predictPC) && (io_output_payload_branchResult_branchResult && io_input_payload_branchInfo_predictResult)) || (io_output_payload_branchResult_branchResult ^ io_input_payload_branchInfo_predictResult));
  always @(*) begin
    case(io_input_payload_uop_bruOp)
      BRUOp_add : begin
        io_output_payload_branchResult_branchResult = 1'b1;
      end
      BRUOp_cadd : begin
        io_output_payload_branchResult_branchResult = io_output_payload_data[0];
      end
      BRUOp_ncadd : begin
        io_output_payload_branchResult_branchResult = io_output_payload_data[0];
      end
      default : begin
        io_output_payload_branchResult_branchResult = 1'b0;
      end
    endcase
  end


endmodule

module ALU (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [31:0]   io_input_payload_src1,
  input  wire [31:0]   io_input_payload_src2,
  input  wire [31:0]   io_input_payload_src3,
  input  wire [31:0]   io_input_payload_src4,
  input  wire [4:0]    io_input_payload_robIdx,
  input  wire [31:0]   io_input_payload_branchInfo_predictPC,
  input  wire          io_input_payload_branchInfo_predictResult,
  input  wire          io_input_payload_exceptionInfo_exception,
  input  wire [5:0]    io_input_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_input_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_payload_pc,
  input  wire [5:0]    io_input_payload_prd,
  input  wire [3:0]    io_input_payload_uop_aluOp,
  input  wire [1:0]    io_input_payload_uop_bruOp,
  input  wire [1:0]    io_input_payload_uop_cruOp,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [4:0]    io_output_payload_robIdx,
  output reg  [31:0]   io_output_payload_data,
  output wire [5:0]    io_output_payload_prd,
  output wire [31:0]   io_output_payload_branchResult_targetPC,
  output reg           io_output_payload_branchResult_branchResult,
  output wire          io_output_payload_branchResult_predictFail,
  output wire          io_output_payload_exceptionInfo_exception,
  output wire [5:0]    io_output_payload_exceptionInfo_eCode,
  output wire [0:0]    io_output_payload_exceptionInfo_eSubCode,
  output wire          io_forward_valid,
  output wire [5:0]    io_forward_payload_idx,
  output wire [31:0]   io_forward_payload_payload,
  output wire          io_wakeOut_valid,
  output wire [5:0]    io_wakeOut_payload,
  output reg  [31:0]   io_csrWrite_value,
  output wire [13:0]   io_csrWrite_address,
  output reg           io_csrWrite_wen
);
  localparam ALUOp_add = 4'd0;
  localparam ALUOp_sub = 4'd1;
  localparam ALUOp_slt = 4'd2;
  localparam ALUOp_sltu = 4'd3;
  localparam ALUOp_eq = 4'd4;
  localparam ALUOp_nor_1 = 4'd5;
  localparam ALUOp_and_1 = 4'd6;
  localparam ALUOp_or_1 = 4'd7;
  localparam ALUOp_xor_1 = 4'd8;
  localparam ALUOp_sll_1 = 4'd9;
  localparam ALUOp_srl_1 = 4'd10;
  localparam ALUOp_sra_1 = 4'd11;
  localparam ALUOp_passa = 4'd12;
  localparam ALUOp_passb = 4'd13;
  localparam BRUOp_nop = 2'd0;
  localparam BRUOp_add = 2'd1;
  localparam BRUOp_cadd = 2'd2;
  localparam BRUOp_ncadd = 2'd3;
  localparam CRUOp_nop = 2'd0;
  localparam CRUOp_pass = 2'd1;
  localparam CRUOp_mask = 2'd2;

  wire       [31:0]   _zz_slt;
  wire       [31:0]   _zz_slt_1;
  wire       [31:0]   _zz_sra_1;
  wire       [31:0]   _zz_sra_1_1;
  wire       [31:0]   _zz_io_csrWrite_address;
  wire       [31:0]   add;
  wire       [31:0]   sub;
  wire       [0:0]    slt;
  wire       [0:0]    sltu;
  wire       [0:0]    eq;
  wire       [31:0]   nor_1;
  wire       [31:0]   and_1;
  wire       [31:0]   or_1;
  wire       [31:0]   xor_1;
  wire       [31:0]   sll_1;
  wire       [31:0]   srl_1;
  wire       [31:0]   sra_1;
  `ifndef SYNTHESIS
  reg [39:0] io_input_payload_uop_aluOp_string;
  reg [39:0] io_input_payload_uop_bruOp_string;
  reg [31:0] io_input_payload_uop_cruOp_string;
  `endif


  assign _zz_slt = io_input_payload_src1;
  assign _zz_slt_1 = io_input_payload_src2;
  assign _zz_sra_1 = ($signed(_zz_sra_1_1) >>> io_input_payload_src2[4 : 0]);
  assign _zz_sra_1_1 = io_input_payload_src1;
  assign _zz_io_csrWrite_address = io_input_payload_src2;
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_uop_aluOp)
      ALUOp_add : io_input_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_input_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_input_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_input_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_input_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_input_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_input_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_input_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_input_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_input_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_input_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_input_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_input_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_input_payload_uop_aluOp_string = "passb";
      default : io_input_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_input_payload_uop_bruOp)
      BRUOp_nop : io_input_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_input_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_input_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_input_payload_uop_bruOp_string = "ncadd";
      default : io_input_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_input_payload_uop_cruOp)
      CRUOp_nop : io_input_payload_uop_cruOp_string = "nop ";
      CRUOp_pass : io_input_payload_uop_cruOp_string = "pass";
      CRUOp_mask : io_input_payload_uop_cruOp_string = "mask";
      default : io_input_payload_uop_cruOp_string = "????";
    endcase
  end
  `endif

  assign io_input_ready = io_output_ready;
  assign io_output_valid = io_input_valid;
  assign io_output_payload_robIdx = io_input_payload_robIdx;
  assign io_output_payload_prd = io_input_payload_prd;
  assign io_output_payload_exceptionInfo_exception = io_input_payload_exceptionInfo_exception;
  assign io_output_payload_exceptionInfo_eCode = io_input_payload_exceptionInfo_eCode;
  assign io_output_payload_exceptionInfo_eSubCode = io_input_payload_exceptionInfo_eSubCode;
  assign io_forward_valid = (io_input_valid && (io_input_payload_prd != 6'h00));
  assign io_forward_payload_idx = io_input_payload_prd;
  assign io_forward_payload_payload = io_output_payload_data;
  assign io_wakeOut_valid = io_input_valid;
  assign io_wakeOut_payload = io_input_payload_prd;
  assign add = (io_input_payload_src1 + io_input_payload_src2);
  assign sub = (io_input_payload_src1 - io_input_payload_src2);
  assign slt = ($signed(_zz_slt) < $signed(_zz_slt_1));
  assign sltu = (io_input_payload_src1 < io_input_payload_src2);
  assign eq = (io_input_payload_src1 == io_input_payload_src2);
  assign nor_1 = (~ (io_input_payload_src1 | io_input_payload_src2));
  assign and_1 = (io_input_payload_src1 & io_input_payload_src2);
  assign or_1 = (io_input_payload_src1 | io_input_payload_src2);
  assign xor_1 = (io_input_payload_src1 ^ io_input_payload_src2);
  assign sll_1 = (io_input_payload_src1 <<< io_input_payload_src2[4 : 0]);
  assign srl_1 = (io_input_payload_src1 >>> io_input_payload_src2[4 : 0]);
  assign sra_1 = _zz_sra_1;
  always @(*) begin
    case(io_input_payload_uop_aluOp)
      ALUOp_add : begin
        io_output_payload_data = add;
      end
      ALUOp_sub : begin
        io_output_payload_data = sub;
      end
      ALUOp_slt : begin
        io_output_payload_data = {31'd0, slt};
      end
      ALUOp_sltu : begin
        io_output_payload_data = {31'd0, sltu};
      end
      ALUOp_eq : begin
        io_output_payload_data = {31'd0, eq};
      end
      ALUOp_nor_1 : begin
        io_output_payload_data = nor_1;
      end
      ALUOp_and_1 : begin
        io_output_payload_data = and_1;
      end
      ALUOp_or_1 : begin
        io_output_payload_data = or_1;
      end
      ALUOp_xor_1 : begin
        io_output_payload_data = xor_1;
      end
      ALUOp_sll_1 : begin
        io_output_payload_data = sll_1;
      end
      ALUOp_srl_1 : begin
        io_output_payload_data = srl_1;
      end
      ALUOp_sra_1 : begin
        io_output_payload_data = sra_1;
      end
      ALUOp_passa : begin
        io_output_payload_data = io_input_payload_src1;
      end
      default : begin
        io_output_payload_data = io_input_payload_src2;
      end
    endcase
  end

  assign io_output_payload_branchResult_targetPC = (io_input_payload_src3 + io_input_payload_src4);
  assign io_output_payload_branchResult_predictFail = (((io_output_payload_branchResult_targetPC != io_input_payload_branchInfo_predictPC) && (io_output_payload_branchResult_branchResult && io_input_payload_branchInfo_predictResult)) || (io_output_payload_branchResult_branchResult ^ io_input_payload_branchInfo_predictResult));
  always @(*) begin
    case(io_input_payload_uop_bruOp)
      BRUOp_add : begin
        io_output_payload_branchResult_branchResult = 1'b1;
      end
      BRUOp_cadd : begin
        io_output_payload_branchResult_branchResult = io_output_payload_data[0];
      end
      BRUOp_ncadd : begin
        io_output_payload_branchResult_branchResult = io_output_payload_data[0];
      end
      default : begin
        io_output_payload_branchResult_branchResult = 1'b0;
      end
    endcase
  end

  assign io_csrWrite_address = _zz_io_csrWrite_address[13:0];
  always @(*) begin
    io_csrWrite_value = io_input_payload_src4;
    case(io_input_payload_uop_cruOp)
      CRUOp_pass : begin
        io_csrWrite_value = io_input_payload_src4;
      end
      CRUOp_mask : begin
        io_csrWrite_value = ((io_input_payload_src4 & io_input_payload_src3) | (io_input_payload_src1 & (~ io_input_payload_src3)));
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_csrWrite_wen = 1'b0;
    case(io_input_payload_uop_cruOp)
      CRUOp_pass : begin
        io_csrWrite_wen = 1'b1;
      end
      CRUOp_mask : begin
        io_csrWrite_wen = 1'b1;
      end
      default : begin
      end
    endcase
  end


endmodule

module ReadOperandLogic_4 (
  input  wire          io_cmd_valid,
  output wire          io_cmd_ready,
  input  wire [4:0]    io_cmd_payload_robIdx,
  input  wire [31:0]   io_cmd_payload_branchResult_targetPC,
  input  wire          io_cmd_payload_branchResult_branchResult,
  input  wire          io_cmd_payload_branchResult_predictFail,
  input  wire          io_cmd_payload_exceptionInfo_exception,
  input  wire [5:0]    io_cmd_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_cmd_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_cmd_payload_pc,
  input  wire [5:0]    io_cmd_payload_prd,
  input  wire [5:0]    io_cmd_payload_psrc_0,
  input  wire [5:0]    io_cmd_payload_psrc_1,
  input  wire [31:0]   io_cmd_payload_imm,
  input  wire [3:0]    io_cmd_payload_uop_lsuOp,
  input  wire [4:0]    io_cmd_payload_uop_lsuCoOp,
  input  wire [0:0]    io_cmd_payload_roop_lsuROOp,
  output wire          io_toFU_valid,
  input  wire          io_toFU_ready,
  output wire [31:0]   io_toFU_payload_src1,
  output reg  [31:0]   io_toFU_payload_src2,
  output wire [31:0]   io_toFU_payload_src3,
  output wire [4:0]    io_toFU_payload_robIdx,
  output wire [31:0]   io_toFU_payload_branchResult_targetPC,
  output wire          io_toFU_payload_branchResult_branchResult,
  output wire          io_toFU_payload_branchResult_predictFail,
  output wire          io_toFU_payload_exceptionInfo_exception,
  output wire [5:0]    io_toFU_payload_exceptionInfo_eCode,
  output wire [0:0]    io_toFU_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_toFU_payload_pc,
  output wire [5:0]    io_toFU_payload_prd,
  output wire [3:0]    io_toFU_payload_uop_lsuOp,
  output wire [4:0]    io_toFU_payload_uop_lsuCoOp,
  input  wire          io_forward_0_valid,
  input  wire [5:0]    io_forward_0_payload_idx,
  input  wire [31:0]   io_forward_0_payload_payload,
  input  wire          io_forward_1_valid,
  input  wire [5:0]    io_forward_1_payload_idx,
  input  wire [31:0]   io_forward_1_payload_payload,
  input  wire          io_forward_2_valid,
  input  wire [5:0]    io_forward_2_payload_idx,
  input  wire [31:0]   io_forward_2_payload_payload,
  input  wire          io_forward_3_valid,
  input  wire [5:0]    io_forward_3_payload_idx,
  input  wire [31:0]   io_forward_3_payload_payload,
  input  wire          io_forward_4_valid,
  input  wire [5:0]    io_forward_4_payload_idx,
  input  wire [31:0]   io_forward_4_payload_payload,
  input  wire          io_forward_5_valid,
  input  wire [5:0]    io_forward_5_payload_idx,
  input  wire [31:0]   io_forward_5_payload_payload,
  input  wire          io_forward_6_valid,
  input  wire [5:0]    io_forward_6_payload_idx,
  input  wire [31:0]   io_forward_6_payload_payload,
  output wire [5:0]    io_prf_0_idx,
  input  wire [31:0]   io_prf_0_data,
  output wire [5:0]    io_prf_1_idx,
  input  wire [31:0]   io_prf_1_data,
  input  wire          io_interrupt
);
  localparam LSUOp_cacop = 4'd0;
  localparam LSUOp_tlbsrch = 4'd1;
  localparam LSUOp_tlbrd = 4'd2;
  localparam LSUOp_tlbwr = 4'd3;
  localparam LSUOp_tlbfill = 4'd4;
  localparam LSUOp_invtlb = 4'd5;
  localparam LSUOp_ll = 4'd6;
  localparam LSUOp_sc = 4'd7;
  localparam LSUOp_ld = 4'd8;
  localparam LSUOp_ldu = 4'd9;
  localparam LSUOp_st = 4'd10;
  localparam LSUOp_preld = 4'd11;
  localparam LSUOp_dbar = 4'd12;
  localparam LSUOp_ibar = 4'd13;
  localparam LSUROOp_reg_1 = 1'd0;
  localparam LSUROOp_regimm = 1'd1;

  wire                interruptInfo_exception;
  wire       [5:0]    interruptInfo_eCode;
  wire       [0:0]    interruptInfo_eSubCode;
  reg        [31:0]   reg1;
  wire                when_ReadOperand_l49;
  wire                when_ReadOperand_l49_1;
  wire                when_ReadOperand_l49_2;
  wire                when_ReadOperand_l49_3;
  wire                when_ReadOperand_l49_4;
  wire                when_ReadOperand_l49_5;
  wire                when_ReadOperand_l49_6;
  reg        [31:0]   reg2;
  wire                when_ReadOperand_l59;
  wire                when_ReadOperand_l59_1;
  wire                when_ReadOperand_l59_2;
  wire                when_ReadOperand_l59_3;
  wire                when_ReadOperand_l59_4;
  wire                when_ReadOperand_l59_5;
  wire                when_ReadOperand_l59_6;
  wire       [31:0]   csr_1;
  `ifndef SYNTHESIS
  reg [55:0] io_cmd_payload_uop_lsuOp_string;
  reg [47:0] io_cmd_payload_roop_lsuROOp_string;
  reg [55:0] io_toFU_payload_uop_lsuOp_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(io_cmd_payload_uop_lsuOp)
      LSUOp_cacop : io_cmd_payload_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : io_cmd_payload_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : io_cmd_payload_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : io_cmd_payload_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : io_cmd_payload_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : io_cmd_payload_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : io_cmd_payload_uop_lsuOp_string = "ll     ";
      LSUOp_sc : io_cmd_payload_uop_lsuOp_string = "sc     ";
      LSUOp_ld : io_cmd_payload_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : io_cmd_payload_uop_lsuOp_string = "ldu    ";
      LSUOp_st : io_cmd_payload_uop_lsuOp_string = "st     ";
      LSUOp_preld : io_cmd_payload_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : io_cmd_payload_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : io_cmd_payload_uop_lsuOp_string = "ibar   ";
      default : io_cmd_payload_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_cmd_payload_roop_lsuROOp)
      LSUROOp_reg_1 : io_cmd_payload_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : io_cmd_payload_roop_lsuROOp_string = "regimm";
      default : io_cmd_payload_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_toFU_payload_uop_lsuOp)
      LSUOp_cacop : io_toFU_payload_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : io_toFU_payload_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : io_toFU_payload_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : io_toFU_payload_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : io_toFU_payload_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : io_toFU_payload_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : io_toFU_payload_uop_lsuOp_string = "ll     ";
      LSUOp_sc : io_toFU_payload_uop_lsuOp_string = "sc     ";
      LSUOp_ld : io_toFU_payload_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : io_toFU_payload_uop_lsuOp_string = "ldu    ";
      LSUOp_st : io_toFU_payload_uop_lsuOp_string = "st     ";
      LSUOp_preld : io_toFU_payload_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : io_toFU_payload_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : io_toFU_payload_uop_lsuOp_string = "ibar   ";
      default : io_toFU_payload_uop_lsuOp_string = "???????";
    endcase
  end
  `endif

  assign io_toFU_payload_robIdx = io_cmd_payload_robIdx;
  assign io_toFU_payload_branchResult_targetPC = io_cmd_payload_branchResult_targetPC;
  assign io_toFU_payload_branchResult_branchResult = io_cmd_payload_branchResult_branchResult;
  assign io_toFU_payload_branchResult_predictFail = io_cmd_payload_branchResult_predictFail;
  assign interruptInfo_exception = 1'b1;
  assign interruptInfo_eCode = 6'h00;
  assign interruptInfo_eSubCode = 1'b0;
  assign io_toFU_payload_exceptionInfo_exception = (io_interrupt ? interruptInfo_exception : io_cmd_payload_exceptionInfo_exception);
  assign io_toFU_payload_exceptionInfo_eCode = (io_interrupt ? interruptInfo_eCode : io_cmd_payload_exceptionInfo_eCode);
  assign io_toFU_payload_exceptionInfo_eSubCode = (io_interrupt ? interruptInfo_eSubCode : io_cmd_payload_exceptionInfo_eSubCode);
  assign io_toFU_payload_pc = io_cmd_payload_pc;
  assign io_toFU_payload_prd = io_cmd_payload_prd;
  assign io_toFU_payload_uop_lsuOp = io_cmd_payload_uop_lsuOp;
  assign io_toFU_payload_uop_lsuCoOp = io_cmd_payload_uop_lsuCoOp;
  assign io_toFU_valid = io_cmd_valid;
  assign io_cmd_ready = io_toFU_ready;
  assign io_prf_0_idx = io_cmd_payload_psrc_0;
  always @(*) begin
    reg1 = io_prf_0_data;
    if(when_ReadOperand_l49) begin
      reg1 = io_forward_0_payload_payload;
    end
    if(when_ReadOperand_l49_1) begin
      reg1 = io_forward_1_payload_payload;
    end
    if(when_ReadOperand_l49_2) begin
      reg1 = io_forward_2_payload_payload;
    end
    if(when_ReadOperand_l49_3) begin
      reg1 = io_forward_3_payload_payload;
    end
    if(when_ReadOperand_l49_4) begin
      reg1 = io_forward_4_payload_payload;
    end
    if(when_ReadOperand_l49_5) begin
      reg1 = io_forward_5_payload_payload;
    end
    if(when_ReadOperand_l49_6) begin
      reg1 = io_forward_6_payload_payload;
    end
  end

  assign when_ReadOperand_l49 = ((io_forward_0_payload_idx == io_cmd_payload_psrc_0) && io_forward_0_valid);
  assign when_ReadOperand_l49_1 = ((io_forward_1_payload_idx == io_cmd_payload_psrc_0) && io_forward_1_valid);
  assign when_ReadOperand_l49_2 = ((io_forward_2_payload_idx == io_cmd_payload_psrc_0) && io_forward_2_valid);
  assign when_ReadOperand_l49_3 = ((io_forward_3_payload_idx == io_cmd_payload_psrc_0) && io_forward_3_valid);
  assign when_ReadOperand_l49_4 = ((io_forward_4_payload_idx == io_cmd_payload_psrc_0) && io_forward_4_valid);
  assign when_ReadOperand_l49_5 = ((io_forward_5_payload_idx == io_cmd_payload_psrc_0) && io_forward_5_valid);
  assign when_ReadOperand_l49_6 = ((io_forward_6_payload_idx == io_cmd_payload_psrc_0) && io_forward_6_valid);
  assign io_prf_1_idx = io_cmd_payload_psrc_1;
  always @(*) begin
    reg2 = io_prf_1_data;
    if(when_ReadOperand_l59) begin
      reg2 = io_forward_0_payload_payload;
    end
    if(when_ReadOperand_l59_1) begin
      reg2 = io_forward_1_payload_payload;
    end
    if(when_ReadOperand_l59_2) begin
      reg2 = io_forward_2_payload_payload;
    end
    if(when_ReadOperand_l59_3) begin
      reg2 = io_forward_3_payload_payload;
    end
    if(when_ReadOperand_l59_4) begin
      reg2 = io_forward_4_payload_payload;
    end
    if(when_ReadOperand_l59_5) begin
      reg2 = io_forward_5_payload_payload;
    end
    if(when_ReadOperand_l59_6) begin
      reg2 = io_forward_6_payload_payload;
    end
  end

  assign when_ReadOperand_l59 = ((io_forward_0_payload_idx == io_cmd_payload_psrc_1) && io_forward_0_valid);
  assign when_ReadOperand_l59_1 = ((io_forward_1_payload_idx == io_cmd_payload_psrc_1) && io_forward_1_valid);
  assign when_ReadOperand_l59_2 = ((io_forward_2_payload_idx == io_cmd_payload_psrc_1) && io_forward_2_valid);
  assign when_ReadOperand_l59_3 = ((io_forward_3_payload_idx == io_cmd_payload_psrc_1) && io_forward_3_valid);
  assign when_ReadOperand_l59_4 = ((io_forward_4_payload_idx == io_cmd_payload_psrc_1) && io_forward_4_valid);
  assign when_ReadOperand_l59_5 = ((io_forward_5_payload_idx == io_cmd_payload_psrc_1) && io_forward_5_valid);
  assign when_ReadOperand_l59_6 = ((io_forward_6_payload_idx == io_cmd_payload_psrc_1) && io_forward_6_valid);
  assign io_toFU_payload_src1 = reg1;
  assign io_toFU_payload_src3 = reg2;
  always @(*) begin
    case(io_cmd_payload_roop_lsuROOp)
      LSUROOp_reg_1 : begin
        io_toFU_payload_src2 = reg2;
      end
      default : begin
        io_toFU_payload_src2 = io_cmd_payload_imm;
      end
    endcase
  end


endmodule

module ReadOperandLogic_3 (
  input  wire          io_cmd_valid,
  output wire          io_cmd_ready,
  input  wire [4:0]    io_cmd_payload_robIdx,
  input  wire [31:0]   io_cmd_payload_branchResult_targetPC,
  input  wire          io_cmd_payload_branchResult_branchResult,
  input  wire          io_cmd_payload_branchResult_predictFail,
  input  wire          io_cmd_payload_exceptionInfo_exception,
  input  wire [5:0]    io_cmd_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_cmd_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_cmd_payload_pc,
  input  wire [5:0]    io_cmd_payload_prd,
  input  wire [5:0]    io_cmd_payload_psrc_0,
  input  wire [5:0]    io_cmd_payload_psrc_1,
  input  wire [31:0]   io_cmd_payload_imm,
  input  wire [1:0]    io_cmd_payload_uop_divuOp,
  output wire          io_toFU_valid,
  input  wire          io_toFU_ready,
  output wire [31:0]   io_toFU_payload_src1,
  output wire [31:0]   io_toFU_payload_src2,
  output wire [4:0]    io_toFU_payload_robIdx,
  output wire [31:0]   io_toFU_payload_branchResult_targetPC,
  output wire          io_toFU_payload_branchResult_branchResult,
  output wire          io_toFU_payload_branchResult_predictFail,
  output wire          io_toFU_payload_exceptionInfo_exception,
  output wire [5:0]    io_toFU_payload_exceptionInfo_eCode,
  output wire [0:0]    io_toFU_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_toFU_payload_pc,
  output wire [5:0]    io_toFU_payload_prd,
  output wire [1:0]    io_toFU_payload_uop_divuOp,
  output wire [5:0]    io_prf_0_idx,
  input  wire [31:0]   io_prf_0_data,
  output wire [5:0]    io_prf_1_idx,
  input  wire [31:0]   io_prf_1_data,
  input  wire          io_interrupt
);
  localparam DIVUOp_div = 2'd0;
  localparam DIVUOp_divu = 2'd1;
  localparam DIVUOp_mod_1 = 2'd2;
  localparam DIVUOp_modu = 2'd3;

  wire                interruptInfo_exception;
  wire       [5:0]    interruptInfo_eCode;
  wire       [0:0]    interruptInfo_eSubCode;
  wire       [31:0]   reg1;
  wire       [31:0]   reg2;
  wire       [31:0]   csr_1;
  `ifndef SYNTHESIS
  reg [39:0] io_cmd_payload_uop_divuOp_string;
  reg [39:0] io_toFU_payload_uop_divuOp_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(io_cmd_payload_uop_divuOp)
      DIVUOp_div : io_cmd_payload_uop_divuOp_string = "div  ";
      DIVUOp_divu : io_cmd_payload_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : io_cmd_payload_uop_divuOp_string = "mod_1";
      DIVUOp_modu : io_cmd_payload_uop_divuOp_string = "modu ";
      default : io_cmd_payload_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_toFU_payload_uop_divuOp)
      DIVUOp_div : io_toFU_payload_uop_divuOp_string = "div  ";
      DIVUOp_divu : io_toFU_payload_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : io_toFU_payload_uop_divuOp_string = "mod_1";
      DIVUOp_modu : io_toFU_payload_uop_divuOp_string = "modu ";
      default : io_toFU_payload_uop_divuOp_string = "?????";
    endcase
  end
  `endif

  assign io_toFU_payload_robIdx = io_cmd_payload_robIdx;
  assign io_toFU_payload_branchResult_targetPC = io_cmd_payload_branchResult_targetPC;
  assign io_toFU_payload_branchResult_branchResult = io_cmd_payload_branchResult_branchResult;
  assign io_toFU_payload_branchResult_predictFail = io_cmd_payload_branchResult_predictFail;
  assign interruptInfo_exception = 1'b1;
  assign interruptInfo_eCode = 6'h00;
  assign interruptInfo_eSubCode = 1'b0;
  assign io_toFU_payload_exceptionInfo_exception = (io_interrupt ? interruptInfo_exception : io_cmd_payload_exceptionInfo_exception);
  assign io_toFU_payload_exceptionInfo_eCode = (io_interrupt ? interruptInfo_eCode : io_cmd_payload_exceptionInfo_eCode);
  assign io_toFU_payload_exceptionInfo_eSubCode = (io_interrupt ? interruptInfo_eSubCode : io_cmd_payload_exceptionInfo_eSubCode);
  assign io_toFU_payload_pc = io_cmd_payload_pc;
  assign io_toFU_payload_prd = io_cmd_payload_prd;
  assign io_toFU_payload_uop_divuOp = io_cmd_payload_uop_divuOp;
  assign io_toFU_valid = io_cmd_valid;
  assign io_cmd_ready = io_toFU_ready;
  assign io_prf_0_idx = io_cmd_payload_psrc_0;
  assign reg1 = io_prf_0_data;
  assign io_prf_1_idx = io_cmd_payload_psrc_1;
  assign reg2 = io_prf_1_data;
  assign io_toFU_payload_src1 = reg1;
  assign io_toFU_payload_src2 = reg2;

endmodule

module ReadOperandLogic_2 (
  input  wire          io_cmd_valid,
  output wire          io_cmd_ready,
  input  wire [4:0]    io_cmd_payload_robIdx,
  input  wire [31:0]   io_cmd_payload_branchResult_targetPC,
  input  wire          io_cmd_payload_branchResult_branchResult,
  input  wire          io_cmd_payload_branchResult_predictFail,
  input  wire          io_cmd_payload_exceptionInfo_exception,
  input  wire [5:0]    io_cmd_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_cmd_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_cmd_payload_pc,
  input  wire [5:0]    io_cmd_payload_prd,
  input  wire [5:0]    io_cmd_payload_psrc_0,
  input  wire [5:0]    io_cmd_payload_psrc_1,
  input  wire [31:0]   io_cmd_payload_imm,
  input  wire [1:0]    io_cmd_payload_uop_muluOp,
  output wire          io_toFU_valid,
  input  wire          io_toFU_ready,
  output wire [31:0]   io_toFU_payload_src1,
  output wire [31:0]   io_toFU_payload_src2,
  output wire [4:0]    io_toFU_payload_robIdx,
  output wire [31:0]   io_toFU_payload_branchResult_targetPC,
  output wire          io_toFU_payload_branchResult_branchResult,
  output wire          io_toFU_payload_branchResult_predictFail,
  output wire          io_toFU_payload_exceptionInfo_exception,
  output wire [5:0]    io_toFU_payload_exceptionInfo_eCode,
  output wire [0:0]    io_toFU_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_toFU_payload_pc,
  output wire [5:0]    io_toFU_payload_prd,
  output wire [1:0]    io_toFU_payload_uop_muluOp,
  input  wire          io_forward_0_valid,
  input  wire [5:0]    io_forward_0_payload_idx,
  input  wire [31:0]   io_forward_0_payload_payload,
  output wire [5:0]    io_prf_0_idx,
  input  wire [31:0]   io_prf_0_data,
  output wire [5:0]    io_prf_1_idx,
  input  wire [31:0]   io_prf_1_data,
  input  wire          io_interrupt
);
  localparam MULUOp_mullo = 2'd0;
  localparam MULUOp_mulhi = 2'd1;
  localparam MULUOp_mulhiu = 2'd2;

  wire                interruptInfo_exception;
  wire       [5:0]    interruptInfo_eCode;
  wire       [0:0]    interruptInfo_eSubCode;
  reg        [31:0]   reg1;
  wire                when_ReadOperand_l49;
  reg        [31:0]   reg2;
  wire                when_ReadOperand_l59;
  wire       [31:0]   csr_1;
  `ifndef SYNTHESIS
  reg [47:0] io_cmd_payload_uop_muluOp_string;
  reg [47:0] io_toFU_payload_uop_muluOp_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(io_cmd_payload_uop_muluOp)
      MULUOp_mullo : io_cmd_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : io_cmd_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : io_cmd_payload_uop_muluOp_string = "mulhiu";
      default : io_cmd_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_toFU_payload_uop_muluOp)
      MULUOp_mullo : io_toFU_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : io_toFU_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : io_toFU_payload_uop_muluOp_string = "mulhiu";
      default : io_toFU_payload_uop_muluOp_string = "??????";
    endcase
  end
  `endif

  assign io_toFU_payload_robIdx = io_cmd_payload_robIdx;
  assign io_toFU_payload_branchResult_targetPC = io_cmd_payload_branchResult_targetPC;
  assign io_toFU_payload_branchResult_branchResult = io_cmd_payload_branchResult_branchResult;
  assign io_toFU_payload_branchResult_predictFail = io_cmd_payload_branchResult_predictFail;
  assign interruptInfo_exception = 1'b1;
  assign interruptInfo_eCode = 6'h00;
  assign interruptInfo_eSubCode = 1'b0;
  assign io_toFU_payload_exceptionInfo_exception = (io_interrupt ? interruptInfo_exception : io_cmd_payload_exceptionInfo_exception);
  assign io_toFU_payload_exceptionInfo_eCode = (io_interrupt ? interruptInfo_eCode : io_cmd_payload_exceptionInfo_eCode);
  assign io_toFU_payload_exceptionInfo_eSubCode = (io_interrupt ? interruptInfo_eSubCode : io_cmd_payload_exceptionInfo_eSubCode);
  assign io_toFU_payload_pc = io_cmd_payload_pc;
  assign io_toFU_payload_prd = io_cmd_payload_prd;
  assign io_toFU_payload_uop_muluOp = io_cmd_payload_uop_muluOp;
  assign io_toFU_valid = io_cmd_valid;
  assign io_cmd_ready = io_toFU_ready;
  assign io_prf_0_idx = io_cmd_payload_psrc_0;
  always @(*) begin
    reg1 = io_prf_0_data;
    if(when_ReadOperand_l49) begin
      reg1 = io_forward_0_payload_payload;
    end
  end

  assign when_ReadOperand_l49 = ((io_forward_0_payload_idx == io_cmd_payload_psrc_0) && io_forward_0_valid);
  assign io_prf_1_idx = io_cmd_payload_psrc_1;
  always @(*) begin
    reg2 = io_prf_1_data;
    if(when_ReadOperand_l59) begin
      reg2 = io_forward_0_payload_payload;
    end
  end

  assign when_ReadOperand_l59 = ((io_forward_0_payload_idx == io_cmd_payload_psrc_1) && io_forward_0_valid);
  assign io_toFU_payload_src1 = reg1;
  assign io_toFU_payload_src2 = reg2;

endmodule

module ReadOperandLogic_1 (
  input  wire          io_cmd_valid,
  output wire          io_cmd_ready,
  input  wire [4:0]    io_cmd_payload_robIdx,
  input  wire [31:0]   io_cmd_payload_branchInfo_predictPC,
  input  wire          io_cmd_payload_branchInfo_predictResult,
  input  wire          io_cmd_payload_exceptionInfo_exception,
  input  wire [5:0]    io_cmd_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_cmd_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_cmd_payload_pc,
  input  wire [5:0]    io_cmd_payload_prd,
  input  wire [5:0]    io_cmd_payload_psrc_0,
  input  wire [5:0]    io_cmd_payload_psrc_1,
  input  wire [31:0]   io_cmd_payload_imm,
  input  wire [3:0]    io_cmd_payload_uop_aluOp,
  input  wire [1:0]    io_cmd_payload_uop_bruOp,
  input  wire [2:0]    io_cmd_payload_roop_aluROOp,
  input  wire [1:0]    io_cmd_payload_roop_cruROOp,
  output wire          io_toFU_valid,
  input  wire          io_toFU_ready,
  output reg  [31:0]   io_toFU_payload_src1,
  output reg  [31:0]   io_toFU_payload_src2,
  output reg  [31:0]   io_toFU_payload_src3,
  output reg  [31:0]   io_toFU_payload_src4,
  output wire [4:0]    io_toFU_payload_robIdx,
  output wire [31:0]   io_toFU_payload_branchInfo_predictPC,
  output wire          io_toFU_payload_branchInfo_predictResult,
  output wire          io_toFU_payload_exceptionInfo_exception,
  output wire [5:0]    io_toFU_payload_exceptionInfo_eCode,
  output wire [0:0]    io_toFU_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_toFU_payload_pc,
  output wire [5:0]    io_toFU_payload_prd,
  output wire [3:0]    io_toFU_payload_uop_aluOp,
  output wire [1:0]    io_toFU_payload_uop_bruOp,
  input  wire          io_forward_0_valid,
  input  wire [5:0]    io_forward_0_payload_idx,
  input  wire [31:0]   io_forward_0_payload_payload,
  input  wire          io_forward_1_valid,
  input  wire [5:0]    io_forward_1_payload_idx,
  input  wire [31:0]   io_forward_1_payload_payload,
  input  wire          io_forward_2_valid,
  input  wire [5:0]    io_forward_2_payload_idx,
  input  wire [31:0]   io_forward_2_payload_payload,
  input  wire          io_forward_3_valid,
  input  wire [5:0]    io_forward_3_payload_idx,
  input  wire [31:0]   io_forward_3_payload_payload,
  input  wire          io_forward_4_valid,
  input  wire [5:0]    io_forward_4_payload_idx,
  input  wire [31:0]   io_forward_4_payload_payload,
  output wire          io_wakeOut_valid,
  output wire [5:0]    io_wakeOut_payload,
  output wire [5:0]    io_prf_0_idx,
  input  wire [31:0]   io_prf_0_data,
  output wire [5:0]    io_prf_1_idx,
  input  wire [31:0]   io_prf_1_data,
  input  wire [31:0]   io_counter_id,
  input  wire [63:0]   io_counter_value,
  input  wire          io_interrupt
);
  localparam ALUOp_add = 4'd0;
  localparam ALUOp_sub = 4'd1;
  localparam ALUOp_slt = 4'd2;
  localparam ALUOp_sltu = 4'd3;
  localparam ALUOp_eq = 4'd4;
  localparam ALUOp_nor_1 = 4'd5;
  localparam ALUOp_and_1 = 4'd6;
  localparam ALUOp_or_1 = 4'd7;
  localparam ALUOp_xor_1 = 4'd8;
  localparam ALUOp_sll_1 = 4'd9;
  localparam ALUOp_srl_1 = 4'd10;
  localparam ALUOp_sra_1 = 4'd11;
  localparam ALUOp_passa = 4'd12;
  localparam ALUOp_passb = 4'd13;
  localparam BRUOp_nop = 2'd0;
  localparam BRUOp_add = 2'd1;
  localparam BRUOp_cadd = 2'd2;
  localparam BRUOp_ncadd = 2'd3;
  localparam ALUROOp_reg_1 = 3'd0;
  localparam ALUROOp_regimm = 3'd1;
  localparam ALUROOp_pcimm = 3'd2;
  localparam ALUROOp_csr = 3'd3;
  localparam ALUROOp_linkpc = 3'd4;
  localparam ALUROOp_linkreg = 3'd5;
  localparam CRUROOp_id = 2'd0;
  localparam CRUROOp_lo = 2'd1;
  localparam CRUROOp_hi = 2'd2;

  wire       [2:0]    _zz_io_toFU_payload_src2;
  wire       [2:0]    _zz_io_toFU_payload_src2_1;
  wire                interruptInfo_exception;
  wire       [5:0]    interruptInfo_eCode;
  wire       [0:0]    interruptInfo_eSubCode;
  reg        [31:0]   reg1;
  wire                when_ReadOperand_l49;
  wire                when_ReadOperand_l49_1;
  wire                when_ReadOperand_l49_2;
  wire                when_ReadOperand_l49_3;
  wire                when_ReadOperand_l49_4;
  reg        [31:0]   reg2;
  wire                when_ReadOperand_l59;
  wire                when_ReadOperand_l59_1;
  wire                when_ReadOperand_l59_2;
  wire                when_ReadOperand_l59_3;
  wire                when_ReadOperand_l59_4;
  reg        [31:0]   csr_1;
  `ifndef SYNTHESIS
  reg [39:0] io_cmd_payload_uop_aluOp_string;
  reg [39:0] io_cmd_payload_uop_bruOp_string;
  reg [55:0] io_cmd_payload_roop_aluROOp_string;
  reg [15:0] io_cmd_payload_roop_cruROOp_string;
  reg [39:0] io_toFU_payload_uop_aluOp_string;
  reg [39:0] io_toFU_payload_uop_bruOp_string;
  `endif


  assign _zz_io_toFU_payload_src2 = 3'b100;
  assign _zz_io_toFU_payload_src2_1 = 3'b100;
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_cmd_payload_uop_aluOp)
      ALUOp_add : io_cmd_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_cmd_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_cmd_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_cmd_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_cmd_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_cmd_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_cmd_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_cmd_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_cmd_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_cmd_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_cmd_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_cmd_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_cmd_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_cmd_payload_uop_aluOp_string = "passb";
      default : io_cmd_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_cmd_payload_uop_bruOp)
      BRUOp_nop : io_cmd_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_cmd_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_cmd_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_cmd_payload_uop_bruOp_string = "ncadd";
      default : io_cmd_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_cmd_payload_roop_aluROOp)
      ALUROOp_reg_1 : io_cmd_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : io_cmd_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : io_cmd_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : io_cmd_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : io_cmd_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : io_cmd_payload_roop_aluROOp_string = "linkreg";
      default : io_cmd_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_cmd_payload_roop_cruROOp)
      CRUROOp_id : io_cmd_payload_roop_cruROOp_string = "id";
      CRUROOp_lo : io_cmd_payload_roop_cruROOp_string = "lo";
      CRUROOp_hi : io_cmd_payload_roop_cruROOp_string = "hi";
      default : io_cmd_payload_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(io_toFU_payload_uop_aluOp)
      ALUOp_add : io_toFU_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_toFU_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_toFU_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_toFU_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_toFU_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_toFU_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_toFU_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_toFU_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_toFU_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_toFU_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_toFU_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_toFU_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_toFU_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_toFU_payload_uop_aluOp_string = "passb";
      default : io_toFU_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_toFU_payload_uop_bruOp)
      BRUOp_nop : io_toFU_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_toFU_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_toFU_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_toFU_payload_uop_bruOp_string = "ncadd";
      default : io_toFU_payload_uop_bruOp_string = "?????";
    endcase
  end
  `endif

  assign io_toFU_payload_robIdx = io_cmd_payload_robIdx;
  assign io_toFU_payload_branchInfo_predictPC = io_cmd_payload_branchInfo_predictPC;
  assign io_toFU_payload_branchInfo_predictResult = io_cmd_payload_branchInfo_predictResult;
  assign io_wakeOut_valid = io_cmd_valid;
  assign io_wakeOut_payload = io_cmd_payload_prd;
  assign interruptInfo_exception = 1'b1;
  assign interruptInfo_eCode = 6'h00;
  assign interruptInfo_eSubCode = 1'b0;
  assign io_toFU_payload_exceptionInfo_exception = (io_interrupt ? interruptInfo_exception : io_cmd_payload_exceptionInfo_exception);
  assign io_toFU_payload_exceptionInfo_eCode = (io_interrupt ? interruptInfo_eCode : io_cmd_payload_exceptionInfo_eCode);
  assign io_toFU_payload_exceptionInfo_eSubCode = (io_interrupt ? interruptInfo_eSubCode : io_cmd_payload_exceptionInfo_eSubCode);
  assign io_toFU_payload_pc = io_cmd_payload_pc;
  assign io_toFU_payload_prd = io_cmd_payload_prd;
  assign io_toFU_payload_uop_aluOp = io_cmd_payload_uop_aluOp;
  assign io_toFU_payload_uop_bruOp = io_cmd_payload_uop_bruOp;
  assign io_toFU_valid = io_cmd_valid;
  assign io_cmd_ready = io_toFU_ready;
  assign io_prf_0_idx = io_cmd_payload_psrc_0;
  always @(*) begin
    reg1 = io_prf_0_data;
    if(when_ReadOperand_l49) begin
      reg1 = io_forward_0_payload_payload;
    end
    if(when_ReadOperand_l49_1) begin
      reg1 = io_forward_1_payload_payload;
    end
    if(when_ReadOperand_l49_2) begin
      reg1 = io_forward_2_payload_payload;
    end
    if(when_ReadOperand_l49_3) begin
      reg1 = io_forward_3_payload_payload;
    end
    if(when_ReadOperand_l49_4) begin
      reg1 = io_forward_4_payload_payload;
    end
  end

  assign when_ReadOperand_l49 = ((io_forward_0_payload_idx == io_cmd_payload_psrc_0) && io_forward_0_valid);
  assign when_ReadOperand_l49_1 = ((io_forward_1_payload_idx == io_cmd_payload_psrc_0) && io_forward_1_valid);
  assign when_ReadOperand_l49_2 = ((io_forward_2_payload_idx == io_cmd_payload_psrc_0) && io_forward_2_valid);
  assign when_ReadOperand_l49_3 = ((io_forward_3_payload_idx == io_cmd_payload_psrc_0) && io_forward_3_valid);
  assign when_ReadOperand_l49_4 = ((io_forward_4_payload_idx == io_cmd_payload_psrc_0) && io_forward_4_valid);
  assign io_prf_1_idx = io_cmd_payload_psrc_1;
  always @(*) begin
    reg2 = io_prf_1_data;
    if(when_ReadOperand_l59) begin
      reg2 = io_forward_0_payload_payload;
    end
    if(when_ReadOperand_l59_1) begin
      reg2 = io_forward_1_payload_payload;
    end
    if(when_ReadOperand_l59_2) begin
      reg2 = io_forward_2_payload_payload;
    end
    if(when_ReadOperand_l59_3) begin
      reg2 = io_forward_3_payload_payload;
    end
    if(when_ReadOperand_l59_4) begin
      reg2 = io_forward_4_payload_payload;
    end
  end

  assign when_ReadOperand_l59 = ((io_forward_0_payload_idx == io_cmd_payload_psrc_1) && io_forward_0_valid);
  assign when_ReadOperand_l59_1 = ((io_forward_1_payload_idx == io_cmd_payload_psrc_1) && io_forward_1_valid);
  assign when_ReadOperand_l59_2 = ((io_forward_2_payload_idx == io_cmd_payload_psrc_1) && io_forward_2_valid);
  assign when_ReadOperand_l59_3 = ((io_forward_3_payload_idx == io_cmd_payload_psrc_1) && io_forward_3_valid);
  assign when_ReadOperand_l59_4 = ((io_forward_4_payload_idx == io_cmd_payload_psrc_1) && io_forward_4_valid);
  always @(*) begin
    case(io_cmd_payload_roop_cruROOp)
      CRUROOp_id : begin
        csr_1 = io_counter_id;
      end
      CRUROOp_lo : begin
        csr_1 = io_counter_value[31 : 0];
      end
      default : begin
        csr_1 = io_counter_value[63 : 32];
      end
    endcase
  end

  always @(*) begin
    case(io_cmd_payload_roop_aluROOp)
      ALUROOp_reg_1 : begin
        io_toFU_payload_src1 = reg1;
      end
      ALUROOp_regimm : begin
        io_toFU_payload_src1 = reg1;
      end
      ALUROOp_pcimm : begin
        io_toFU_payload_src1 = io_cmd_payload_pc;
      end
      ALUROOp_csr : begin
        io_toFU_payload_src1 = csr_1;
      end
      ALUROOp_linkpc : begin
        io_toFU_payload_src1 = io_cmd_payload_pc;
      end
      default : begin
        io_toFU_payload_src1 = io_cmd_payload_pc;
      end
    endcase
  end

  always @(*) begin
    case(io_cmd_payload_roop_aluROOp)
      ALUROOp_reg_1 : begin
        io_toFU_payload_src2 = reg2;
      end
      ALUROOp_regimm : begin
        io_toFU_payload_src2 = io_cmd_payload_imm;
      end
      ALUROOp_pcimm : begin
        io_toFU_payload_src2 = io_cmd_payload_imm;
      end
      ALUROOp_csr : begin
        io_toFU_payload_src2 = io_cmd_payload_imm;
      end
      ALUROOp_linkpc : begin
        io_toFU_payload_src2 = {29'd0, _zz_io_toFU_payload_src2};
      end
      default : begin
        io_toFU_payload_src2 = {29'd0, _zz_io_toFU_payload_src2_1};
      end
    endcase
  end

  always @(*) begin
    case(io_cmd_payload_roop_aluROOp)
      ALUROOp_reg_1 : begin
        io_toFU_payload_src3 = (io_cmd_payload_imm <<< 2);
      end
      ALUROOp_regimm : begin
        io_toFU_payload_src3 = io_cmd_payload_imm;
      end
      ALUROOp_pcimm : begin
        io_toFU_payload_src3 = io_cmd_payload_imm;
      end
      ALUROOp_csr : begin
        io_toFU_payload_src3 = reg2;
      end
      ALUROOp_linkpc : begin
        io_toFU_payload_src3 = (io_cmd_payload_imm <<< 2);
      end
      default : begin
        io_toFU_payload_src3 = (io_cmd_payload_imm <<< 2);
      end
    endcase
  end

  always @(*) begin
    case(io_cmd_payload_roop_aluROOp)
      ALUROOp_reg_1 : begin
        io_toFU_payload_src4 = io_cmd_payload_pc;
      end
      ALUROOp_regimm : begin
        io_toFU_payload_src4 = io_cmd_payload_pc;
      end
      ALUROOp_pcimm : begin
        io_toFU_payload_src4 = io_cmd_payload_pc;
      end
      ALUROOp_csr : begin
        io_toFU_payload_src4 = reg1;
      end
      ALUROOp_linkpc : begin
        io_toFU_payload_src4 = io_cmd_payload_pc;
      end
      default : begin
        io_toFU_payload_src4 = reg1;
      end
    endcase
  end


endmodule

module ReadOperandLogic (
  input  wire          io_cmd_valid,
  output wire          io_cmd_ready,
  input  wire [4:0]    io_cmd_payload_robIdx,
  input  wire [31:0]   io_cmd_payload_branchInfo_predictPC,
  input  wire          io_cmd_payload_branchInfo_predictResult,
  input  wire          io_cmd_payload_exceptionInfo_exception,
  input  wire [5:0]    io_cmd_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_cmd_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_cmd_payload_pc,
  input  wire [5:0]    io_cmd_payload_prd,
  input  wire [5:0]    io_cmd_payload_psrc_0,
  input  wire [5:0]    io_cmd_payload_psrc_1,
  input  wire [31:0]   io_cmd_payload_imm,
  input  wire [3:0]    io_cmd_payload_uop_aluOp,
  input  wire [1:0]    io_cmd_payload_uop_bruOp,
  input  wire [1:0]    io_cmd_payload_uop_cruOp,
  input  wire [2:0]    io_cmd_payload_roop_aluROOp,
  output wire          io_toFU_valid,
  input  wire          io_toFU_ready,
  output reg  [31:0]   io_toFU_payload_src1,
  output reg  [31:0]   io_toFU_payload_src2,
  output reg  [31:0]   io_toFU_payload_src3,
  output reg  [31:0]   io_toFU_payload_src4,
  output wire [4:0]    io_toFU_payload_robIdx,
  output wire [31:0]   io_toFU_payload_branchInfo_predictPC,
  output wire          io_toFU_payload_branchInfo_predictResult,
  output wire          io_toFU_payload_exceptionInfo_exception,
  output wire [5:0]    io_toFU_payload_exceptionInfo_eCode,
  output wire [0:0]    io_toFU_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_toFU_payload_pc,
  output wire [5:0]    io_toFU_payload_prd,
  output wire [3:0]    io_toFU_payload_uop_aluOp,
  output wire [1:0]    io_toFU_payload_uop_bruOp,
  output wire [1:0]    io_toFU_payload_uop_cruOp,
  input  wire          io_forward_0_valid,
  input  wire [5:0]    io_forward_0_payload_idx,
  input  wire [31:0]   io_forward_0_payload_payload,
  input  wire          io_forward_1_valid,
  input  wire [5:0]    io_forward_1_payload_idx,
  input  wire [31:0]   io_forward_1_payload_payload,
  input  wire          io_forward_2_valid,
  input  wire [5:0]    io_forward_2_payload_idx,
  input  wire [31:0]   io_forward_2_payload_payload,
  input  wire          io_forward_3_valid,
  input  wire [5:0]    io_forward_3_payload_idx,
  input  wire [31:0]   io_forward_3_payload_payload,
  input  wire          io_forward_4_valid,
  input  wire [5:0]    io_forward_4_payload_idx,
  input  wire [31:0]   io_forward_4_payload_payload,
  output wire          io_wakeOut_valid,
  output wire [5:0]    io_wakeOut_payload,
  output wire [5:0]    io_prf_0_idx,
  input  wire [31:0]   io_prf_0_data,
  output wire [5:0]    io_prf_1_idx,
  input  wire [31:0]   io_prf_1_data,
  input  wire [31:0]   io_csr_value,
  output wire [13:0]   io_csr_address,
  input  wire          io_interrupt
);
  localparam ALUOp_add = 4'd0;
  localparam ALUOp_sub = 4'd1;
  localparam ALUOp_slt = 4'd2;
  localparam ALUOp_sltu = 4'd3;
  localparam ALUOp_eq = 4'd4;
  localparam ALUOp_nor_1 = 4'd5;
  localparam ALUOp_and_1 = 4'd6;
  localparam ALUOp_or_1 = 4'd7;
  localparam ALUOp_xor_1 = 4'd8;
  localparam ALUOp_sll_1 = 4'd9;
  localparam ALUOp_srl_1 = 4'd10;
  localparam ALUOp_sra_1 = 4'd11;
  localparam ALUOp_passa = 4'd12;
  localparam ALUOp_passb = 4'd13;
  localparam BRUOp_nop = 2'd0;
  localparam BRUOp_add = 2'd1;
  localparam BRUOp_cadd = 2'd2;
  localparam BRUOp_ncadd = 2'd3;
  localparam CRUOp_nop = 2'd0;
  localparam CRUOp_pass = 2'd1;
  localparam CRUOp_mask = 2'd2;
  localparam ALUROOp_reg_1 = 3'd0;
  localparam ALUROOp_regimm = 3'd1;
  localparam ALUROOp_pcimm = 3'd2;
  localparam ALUROOp_csr = 3'd3;
  localparam ALUROOp_linkpc = 3'd4;
  localparam ALUROOp_linkreg = 3'd5;

  wire       [2:0]    _zz_io_toFU_payload_src2;
  wire       [2:0]    _zz_io_toFU_payload_src2_1;
  wire                interruptInfo_exception;
  wire       [5:0]    interruptInfo_eCode;
  wire       [0:0]    interruptInfo_eSubCode;
  reg        [31:0]   reg1;
  wire                when_ReadOperand_l49;
  wire                when_ReadOperand_l49_1;
  wire                when_ReadOperand_l49_2;
  wire                when_ReadOperand_l49_3;
  wire                when_ReadOperand_l49_4;
  reg        [31:0]   reg2;
  wire                when_ReadOperand_l59;
  wire                when_ReadOperand_l59_1;
  wire                when_ReadOperand_l59_2;
  wire                when_ReadOperand_l59_3;
  wire                when_ReadOperand_l59_4;
  wire       [31:0]   csr_1;
  `ifndef SYNTHESIS
  reg [39:0] io_cmd_payload_uop_aluOp_string;
  reg [39:0] io_cmd_payload_uop_bruOp_string;
  reg [31:0] io_cmd_payload_uop_cruOp_string;
  reg [55:0] io_cmd_payload_roop_aluROOp_string;
  reg [39:0] io_toFU_payload_uop_aluOp_string;
  reg [39:0] io_toFU_payload_uop_bruOp_string;
  reg [31:0] io_toFU_payload_uop_cruOp_string;
  `endif


  assign _zz_io_toFU_payload_src2 = 3'b100;
  assign _zz_io_toFU_payload_src2_1 = 3'b100;
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_cmd_payload_uop_aluOp)
      ALUOp_add : io_cmd_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_cmd_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_cmd_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_cmd_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_cmd_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_cmd_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_cmd_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_cmd_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_cmd_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_cmd_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_cmd_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_cmd_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_cmd_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_cmd_payload_uop_aluOp_string = "passb";
      default : io_cmd_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_cmd_payload_uop_bruOp)
      BRUOp_nop : io_cmd_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_cmd_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_cmd_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_cmd_payload_uop_bruOp_string = "ncadd";
      default : io_cmd_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_cmd_payload_uop_cruOp)
      CRUOp_nop : io_cmd_payload_uop_cruOp_string = "nop ";
      CRUOp_pass : io_cmd_payload_uop_cruOp_string = "pass";
      CRUOp_mask : io_cmd_payload_uop_cruOp_string = "mask";
      default : io_cmd_payload_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(io_cmd_payload_roop_aluROOp)
      ALUROOp_reg_1 : io_cmd_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : io_cmd_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : io_cmd_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : io_cmd_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : io_cmd_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : io_cmd_payload_roop_aluROOp_string = "linkreg";
      default : io_cmd_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_toFU_payload_uop_aluOp)
      ALUOp_add : io_toFU_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_toFU_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_toFU_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_toFU_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_toFU_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_toFU_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_toFU_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_toFU_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_toFU_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_toFU_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_toFU_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_toFU_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_toFU_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_toFU_payload_uop_aluOp_string = "passb";
      default : io_toFU_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_toFU_payload_uop_bruOp)
      BRUOp_nop : io_toFU_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_toFU_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_toFU_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_toFU_payload_uop_bruOp_string = "ncadd";
      default : io_toFU_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_toFU_payload_uop_cruOp)
      CRUOp_nop : io_toFU_payload_uop_cruOp_string = "nop ";
      CRUOp_pass : io_toFU_payload_uop_cruOp_string = "pass";
      CRUOp_mask : io_toFU_payload_uop_cruOp_string = "mask";
      default : io_toFU_payload_uop_cruOp_string = "????";
    endcase
  end
  `endif

  assign io_toFU_payload_robIdx = io_cmd_payload_robIdx;
  assign io_toFU_payload_branchInfo_predictPC = io_cmd_payload_branchInfo_predictPC;
  assign io_toFU_payload_branchInfo_predictResult = io_cmd_payload_branchInfo_predictResult;
  assign io_wakeOut_valid = io_cmd_valid;
  assign io_wakeOut_payload = io_cmd_payload_prd;
  assign interruptInfo_exception = 1'b1;
  assign interruptInfo_eCode = 6'h00;
  assign interruptInfo_eSubCode = 1'b0;
  assign io_toFU_payload_exceptionInfo_exception = (io_interrupt ? interruptInfo_exception : io_cmd_payload_exceptionInfo_exception);
  assign io_toFU_payload_exceptionInfo_eCode = (io_interrupt ? interruptInfo_eCode : io_cmd_payload_exceptionInfo_eCode);
  assign io_toFU_payload_exceptionInfo_eSubCode = (io_interrupt ? interruptInfo_eSubCode : io_cmd_payload_exceptionInfo_eSubCode);
  assign io_toFU_payload_pc = io_cmd_payload_pc;
  assign io_toFU_payload_prd = io_cmd_payload_prd;
  assign io_toFU_payload_uop_aluOp = io_cmd_payload_uop_aluOp;
  assign io_toFU_payload_uop_bruOp = io_cmd_payload_uop_bruOp;
  assign io_toFU_payload_uop_cruOp = io_cmd_payload_uop_cruOp;
  assign io_toFU_valid = io_cmd_valid;
  assign io_cmd_ready = io_toFU_ready;
  assign io_prf_0_idx = io_cmd_payload_psrc_0;
  always @(*) begin
    reg1 = io_prf_0_data;
    if(when_ReadOperand_l49) begin
      reg1 = io_forward_0_payload_payload;
    end
    if(when_ReadOperand_l49_1) begin
      reg1 = io_forward_1_payload_payload;
    end
    if(when_ReadOperand_l49_2) begin
      reg1 = io_forward_2_payload_payload;
    end
    if(when_ReadOperand_l49_3) begin
      reg1 = io_forward_3_payload_payload;
    end
    if(when_ReadOperand_l49_4) begin
      reg1 = io_forward_4_payload_payload;
    end
  end

  assign when_ReadOperand_l49 = ((io_forward_0_payload_idx == io_cmd_payload_psrc_0) && io_forward_0_valid);
  assign when_ReadOperand_l49_1 = ((io_forward_1_payload_idx == io_cmd_payload_psrc_0) && io_forward_1_valid);
  assign when_ReadOperand_l49_2 = ((io_forward_2_payload_idx == io_cmd_payload_psrc_0) && io_forward_2_valid);
  assign when_ReadOperand_l49_3 = ((io_forward_3_payload_idx == io_cmd_payload_psrc_0) && io_forward_3_valid);
  assign when_ReadOperand_l49_4 = ((io_forward_4_payload_idx == io_cmd_payload_psrc_0) && io_forward_4_valid);
  assign io_prf_1_idx = io_cmd_payload_psrc_1;
  always @(*) begin
    reg2 = io_prf_1_data;
    if(when_ReadOperand_l59) begin
      reg2 = io_forward_0_payload_payload;
    end
    if(when_ReadOperand_l59_1) begin
      reg2 = io_forward_1_payload_payload;
    end
    if(when_ReadOperand_l59_2) begin
      reg2 = io_forward_2_payload_payload;
    end
    if(when_ReadOperand_l59_3) begin
      reg2 = io_forward_3_payload_payload;
    end
    if(when_ReadOperand_l59_4) begin
      reg2 = io_forward_4_payload_payload;
    end
  end

  assign when_ReadOperand_l59 = ((io_forward_0_payload_idx == io_cmd_payload_psrc_1) && io_forward_0_valid);
  assign when_ReadOperand_l59_1 = ((io_forward_1_payload_idx == io_cmd_payload_psrc_1) && io_forward_1_valid);
  assign when_ReadOperand_l59_2 = ((io_forward_2_payload_idx == io_cmd_payload_psrc_1) && io_forward_2_valid);
  assign when_ReadOperand_l59_3 = ((io_forward_3_payload_idx == io_cmd_payload_psrc_1) && io_forward_3_valid);
  assign when_ReadOperand_l59_4 = ((io_forward_4_payload_idx == io_cmd_payload_psrc_1) && io_forward_4_valid);
  assign io_csr_address = io_cmd_payload_imm[13 : 0];
  assign csr_1 = io_csr_value;
  always @(*) begin
    case(io_cmd_payload_roop_aluROOp)
      ALUROOp_reg_1 : begin
        io_toFU_payload_src1 = reg1;
      end
      ALUROOp_regimm : begin
        io_toFU_payload_src1 = reg1;
      end
      ALUROOp_pcimm : begin
        io_toFU_payload_src1 = io_cmd_payload_pc;
      end
      ALUROOp_csr : begin
        io_toFU_payload_src1 = csr_1;
      end
      ALUROOp_linkpc : begin
        io_toFU_payload_src1 = io_cmd_payload_pc;
      end
      default : begin
        io_toFU_payload_src1 = io_cmd_payload_pc;
      end
    endcase
  end

  always @(*) begin
    case(io_cmd_payload_roop_aluROOp)
      ALUROOp_reg_1 : begin
        io_toFU_payload_src2 = reg2;
      end
      ALUROOp_regimm : begin
        io_toFU_payload_src2 = io_cmd_payload_imm;
      end
      ALUROOp_pcimm : begin
        io_toFU_payload_src2 = io_cmd_payload_imm;
      end
      ALUROOp_csr : begin
        io_toFU_payload_src2 = io_cmd_payload_imm;
      end
      ALUROOp_linkpc : begin
        io_toFU_payload_src2 = {29'd0, _zz_io_toFU_payload_src2};
      end
      default : begin
        io_toFU_payload_src2 = {29'd0, _zz_io_toFU_payload_src2_1};
      end
    endcase
  end

  always @(*) begin
    case(io_cmd_payload_roop_aluROOp)
      ALUROOp_reg_1 : begin
        io_toFU_payload_src3 = (io_cmd_payload_imm <<< 2);
      end
      ALUROOp_regimm : begin
        io_toFU_payload_src3 = io_cmd_payload_imm;
      end
      ALUROOp_pcimm : begin
        io_toFU_payload_src3 = io_cmd_payload_imm;
      end
      ALUROOp_csr : begin
        io_toFU_payload_src3 = reg2;
      end
      ALUROOp_linkpc : begin
        io_toFU_payload_src3 = (io_cmd_payload_imm <<< 2);
      end
      default : begin
        io_toFU_payload_src3 = (io_cmd_payload_imm <<< 2);
      end
    endcase
  end

  always @(*) begin
    case(io_cmd_payload_roop_aluROOp)
      ALUROOp_reg_1 : begin
        io_toFU_payload_src4 = io_cmd_payload_pc;
      end
      ALUROOp_regimm : begin
        io_toFU_payload_src4 = io_cmd_payload_pc;
      end
      ALUROOp_pcimm : begin
        io_toFU_payload_src4 = io_cmd_payload_pc;
      end
      ALUROOp_csr : begin
        io_toFU_payload_src4 = reg1;
      end
      ALUROOp_linkpc : begin
        io_toFU_payload_src4 = io_cmd_payload_pc;
      end
      default : begin
        io_toFU_payload_src4 = reg1;
      end
    endcase
  end


endmodule

module IssueQueue_4 (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [4:0]    io_input_payload_robIdx,
  input  wire [31:0]   io_input_payload_branchResult_targetPC,
  input  wire          io_input_payload_branchResult_branchResult,
  input  wire          io_input_payload_branchResult_predictFail,
  input  wire          io_input_payload_exceptionInfo_exception,
  input  wire [5:0]    io_input_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_input_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_payload_pc,
  input  wire [5:0]    io_input_payload_prd,
  input  wire [5:0]    io_input_payload_psrc_0,
  input  wire [5:0]    io_input_payload_psrc_1,
  input  wire [31:0]   io_input_payload_imm,
  input  wire [3:0]    io_input_payload_uop_lsuOp,
  input  wire [4:0]    io_input_payload_uop_lsuCoOp,
  input  wire [0:0]    io_input_payload_roop_lsuROOp,
  input  wire          io_input_payload_srcReady_0,
  input  wire          io_input_payload_srcReady_1,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [4:0]    io_output_payload_robIdx,
  output wire [31:0]   io_output_payload_branchResult_targetPC,
  output wire          io_output_payload_branchResult_branchResult,
  output wire          io_output_payload_branchResult_predictFail,
  output wire          io_output_payload_exceptionInfo_exception,
  output wire [5:0]    io_output_payload_exceptionInfo_eCode,
  output wire [0:0]    io_output_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_output_payload_pc,
  output wire [5:0]    io_output_payload_prd,
  output wire [5:0]    io_output_payload_psrc_0,
  output wire [5:0]    io_output_payload_psrc_1,
  output wire [31:0]   io_output_payload_imm,
  output wire [3:0]    io_output_payload_uop_lsuOp,
  output wire [4:0]    io_output_payload_uop_lsuCoOp,
  output wire [0:0]    io_output_payload_roop_lsuROOp,
  input  wire [5:0]    io_writebackSignal_0,
  input  wire [5:0]    io_writebackSignal_1,
  input  wire [5:0]    io_writebackSignal_2,
  input  wire [5:0]    io_writebackSignal_3,
  input  wire [5:0]    io_writebackSignal_4,
  input  wire          io_earlyWakeup_0_valid,
  input  wire [5:0]    io_earlyWakeup_0_payload,
  input  wire          io_earlyWakeup_1_valid,
  input  wire [5:0]    io_earlyWakeup_1_payload,
  input  wire          io_earlyWakeup_2_valid,
  input  wire [5:0]    io_earlyWakeup_2_payload,
  input  wire          io_earlyWakeup_3_valid,
  input  wire [5:0]    io_earlyWakeup_3_payload,
  input  wire          io_earlyWakeup_4_valid,
  input  wire [5:0]    io_earlyWakeup_4_payload,
  input  wire          io_earlyWakeup_5_valid,
  input  wire [5:0]    io_earlyWakeup_5_payload,
  input  wire          io_earlyWakeup_6_valid,
  input  wire [5:0]    io_earlyWakeup_6_payload,
  input  wire          io_earlyWakeup_7_valid,
  input  wire [5:0]    io_earlyWakeup_7_payload,
  input  wire          io_earlyWakeup_8_valid,
  input  wire [5:0]    io_earlyWakeup_8_payload,
  input  wire          io_earlyWakeup_9_valid,
  input  wire [5:0]    io_earlyWakeup_9_payload,
  input  wire          io_earlyWakeup_10_valid,
  input  wire [5:0]    io_earlyWakeup_10_payload,
  input  wire          aclk,
  input  wire          cpuClockingArea_areaFlushReset_newReset
);
  localparam LSUOp_cacop = 4'd0;
  localparam LSUOp_tlbsrch = 4'd1;
  localparam LSUOp_tlbrd = 4'd2;
  localparam LSUOp_tlbwr = 4'd3;
  localparam LSUOp_tlbfill = 4'd4;
  localparam LSUOp_invtlb = 4'd5;
  localparam LSUOp_ll = 4'd6;
  localparam LSUOp_sc = 4'd7;
  localparam LSUOp_ld = 4'd8;
  localparam LSUOp_ldu = 4'd9;
  localparam LSUOp_st = 4'd10;
  localparam LSUOp_preld = 4'd11;
  localparam LSUOp_dbar = 4'd12;
  localparam LSUOp_ibar = 4'd13;
  localparam LSUROOp_reg_1 = 1'd0;
  localparam LSUROOp_regimm = 1'd1;

  wire       [3:0]    _zz_readyToIssue_ohFirst_masked;
  wire       [4:0]    _zz_emptyEntry_ohFirst_masked;
  wire                _zz_appendEntry_srcReady_0;
  wire       [0:0]    _zz_appendEntry_srcReady_0_1;
  wire       [1:0]    _zz_appendEntry_srcReady_0_2;
  wire                _zz_appendEntry_srcReady_0_3;
  wire                _zz_appendEntry_srcReady_0_4;
  wire       [0:0]    _zz_appendEntry_srcReady_0_5;
  wire       [6:0]    _zz_appendEntry_srcReady_0_6;
  wire                _zz_appendEntry_srcReady_0_7;
  wire                _zz_appendEntry_srcReady_0_8;
  wire       [0:0]    _zz_appendEntry_srcReady_0_9;
  wire       [2:0]    _zz_appendEntry_srcReady_0_10;
  wire                _zz_appendEntry_srcReady_1;
  wire       [0:0]    _zz_appendEntry_srcReady_1_1;
  wire       [0:0]    _zz_appendEntry_srcReady_1_2;
  wire                _zz_appendEntry_srcReady_1_3;
  wire                _zz_appendEntry_srcReady_1_4;
  wire       [0:0]    _zz_appendEntry_srcReady_1_5;
  wire       [5:0]    _zz_appendEntry_srcReady_1_6;
  wire                _zz_appendEntry_srcReady_1_7;
  wire                _zz_appendEntry_srcReady_1_8;
  wire       [0:0]    _zz_appendEntry_srcReady_1_9;
  wire       [0:0]    _zz_appendEntry_srcReady_1_10;
  wire                _zz_updatedEntry_0_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_0_2;
  wire                _zz_updatedEntry_0_srcReady_0_3;
  wire                _zz_updatedEntry_0_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_0_5;
  wire       [5:0]    _zz_updatedEntry_0_srcReady_0_6;
  wire                _zz_updatedEntry_0_srcReady_0_7;
  wire                _zz_updatedEntry_0_srcReady_0_8;
  wire                _zz_updatedEntry_0_srcReady_0_9;
  wire                _zz_updatedEntry_0_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_1_2;
  wire                _zz_updatedEntry_0_srcReady_1_3;
  wire                _zz_updatedEntry_0_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_1_5;
  wire       [5:0]    _zz_updatedEntry_0_srcReady_1_6;
  wire                _zz_updatedEntry_0_srcReady_1_7;
  wire                _zz_updatedEntry_0_srcReady_1_8;
  wire                _zz_updatedEntry_0_srcReady_1_9;
  wire                _zz_updatedEntry_1_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_0_2;
  wire                _zz_updatedEntry_1_srcReady_0_3;
  wire                _zz_updatedEntry_1_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_0_5;
  wire       [5:0]    _zz_updatedEntry_1_srcReady_0_6;
  wire                _zz_updatedEntry_1_srcReady_0_7;
  wire                _zz_updatedEntry_1_srcReady_0_8;
  wire                _zz_updatedEntry_1_srcReady_0_9;
  wire                _zz_updatedEntry_1_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_1_2;
  wire                _zz_updatedEntry_1_srcReady_1_3;
  wire                _zz_updatedEntry_1_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_1_5;
  wire       [5:0]    _zz_updatedEntry_1_srcReady_1_6;
  wire                _zz_updatedEntry_1_srcReady_1_7;
  wire                _zz_updatedEntry_1_srcReady_1_8;
  wire                _zz_updatedEntry_1_srcReady_1_9;
  wire                _zz_updatedEntry_2_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_0_2;
  wire                _zz_updatedEntry_2_srcReady_0_3;
  wire                _zz_updatedEntry_2_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_0_5;
  wire       [5:0]    _zz_updatedEntry_2_srcReady_0_6;
  wire                _zz_updatedEntry_2_srcReady_0_7;
  wire                _zz_updatedEntry_2_srcReady_0_8;
  wire                _zz_updatedEntry_2_srcReady_0_9;
  wire                _zz_updatedEntry_2_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_1_2;
  wire                _zz_updatedEntry_2_srcReady_1_3;
  wire                _zz_updatedEntry_2_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_1_5;
  wire       [5:0]    _zz_updatedEntry_2_srcReady_1_6;
  wire                _zz_updatedEntry_2_srcReady_1_7;
  wire                _zz_updatedEntry_2_srcReady_1_8;
  wire                _zz_updatedEntry_2_srcReady_1_9;
  wire                _zz_updatedEntry_3_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_0_2;
  wire                _zz_updatedEntry_3_srcReady_0_3;
  wire                _zz_updatedEntry_3_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_0_5;
  wire       [5:0]    _zz_updatedEntry_3_srcReady_0_6;
  wire                _zz_updatedEntry_3_srcReady_0_7;
  wire                _zz_updatedEntry_3_srcReady_0_8;
  wire                _zz_updatedEntry_3_srcReady_0_9;
  wire                _zz_updatedEntry_3_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_1_2;
  wire                _zz_updatedEntry_3_srcReady_1_3;
  wire                _zz_updatedEntry_3_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_1_5;
  wire       [5:0]    _zz_updatedEntry_3_srcReady_1_6;
  wire                _zz_updatedEntry_3_srcReady_1_7;
  wire                _zz_updatedEntry_3_srcReady_1_8;
  wire                _zz_updatedEntry_3_srcReady_1_9;
  reg                 _zz_issueEntry_valid_4;
  reg        [4:0]    _zz_issueEntry_robIdx;
  reg        [31:0]   _zz_issueEntry_branchResult_targetPC;
  reg                 _zz_issueEntry_branchResult_branchResult;
  reg                 _zz_issueEntry_branchResult_predictFail;
  reg                 _zz_issueEntry_exceptionInfo_exception;
  reg        [5:0]    _zz_issueEntry_exceptionInfo_eCode;
  reg        [0:0]    _zz_issueEntry_exceptionInfo_eSubCode;
  reg        [31:0]   _zz_issueEntry_pc;
  reg        [5:0]    _zz_issueEntry_prd;
  reg        [5:0]    _zz_issueEntry_psrc_0;
  reg        [5:0]    _zz_issueEntry_psrc_1;
  reg        [31:0]   _zz_issueEntry_imm;
  reg        [3:0]    _zz_issueEntry_uop_lsuOp;
  reg        [4:0]    _zz_issueEntry_uop_lsuCoOp;
  reg        [0:0]    _zz_issueEntry_roop_lsuROOp;
  reg                 _zz_issueEntry_srcReady_0;
  reg                 _zz_issueEntry_srcReady_1;
  reg                 queue_0_valid;
  reg        [4:0]    queue_0_robIdx;
  reg        [31:0]   queue_0_branchResult_targetPC;
  reg                 queue_0_branchResult_branchResult;
  reg                 queue_0_branchResult_predictFail;
  reg                 queue_0_exceptionInfo_exception;
  reg        [5:0]    queue_0_exceptionInfo_eCode;
  reg        [0:0]    queue_0_exceptionInfo_eSubCode;
  reg        [31:0]   queue_0_pc;
  reg        [5:0]    queue_0_prd;
  reg        [5:0]    queue_0_psrc_0;
  reg        [5:0]    queue_0_psrc_1;
  reg        [31:0]   queue_0_imm;
  reg        [3:0]    queue_0_uop_lsuOp;
  reg        [4:0]    queue_0_uop_lsuCoOp;
  reg        [0:0]    queue_0_roop_lsuROOp;
  reg                 queue_0_srcReady_0;
  reg                 queue_0_srcReady_1;
  reg                 queue_1_valid;
  reg        [4:0]    queue_1_robIdx;
  reg        [31:0]   queue_1_branchResult_targetPC;
  reg                 queue_1_branchResult_branchResult;
  reg                 queue_1_branchResult_predictFail;
  reg                 queue_1_exceptionInfo_exception;
  reg        [5:0]    queue_1_exceptionInfo_eCode;
  reg        [0:0]    queue_1_exceptionInfo_eSubCode;
  reg        [31:0]   queue_1_pc;
  reg        [5:0]    queue_1_prd;
  reg        [5:0]    queue_1_psrc_0;
  reg        [5:0]    queue_1_psrc_1;
  reg        [31:0]   queue_1_imm;
  reg        [3:0]    queue_1_uop_lsuOp;
  reg        [4:0]    queue_1_uop_lsuCoOp;
  reg        [0:0]    queue_1_roop_lsuROOp;
  reg                 queue_1_srcReady_0;
  reg                 queue_1_srcReady_1;
  reg                 queue_2_valid;
  reg        [4:0]    queue_2_robIdx;
  reg        [31:0]   queue_2_branchResult_targetPC;
  reg                 queue_2_branchResult_branchResult;
  reg                 queue_2_branchResult_predictFail;
  reg                 queue_2_exceptionInfo_exception;
  reg        [5:0]    queue_2_exceptionInfo_eCode;
  reg        [0:0]    queue_2_exceptionInfo_eSubCode;
  reg        [31:0]   queue_2_pc;
  reg        [5:0]    queue_2_prd;
  reg        [5:0]    queue_2_psrc_0;
  reg        [5:0]    queue_2_psrc_1;
  reg        [31:0]   queue_2_imm;
  reg        [3:0]    queue_2_uop_lsuOp;
  reg        [4:0]    queue_2_uop_lsuCoOp;
  reg        [0:0]    queue_2_roop_lsuROOp;
  reg                 queue_2_srcReady_0;
  reg                 queue_2_srcReady_1;
  reg                 queue_3_valid;
  reg        [4:0]    queue_3_robIdx;
  reg        [31:0]   queue_3_branchResult_targetPC;
  reg                 queue_3_branchResult_branchResult;
  reg                 queue_3_branchResult_predictFail;
  reg                 queue_3_exceptionInfo_exception;
  reg        [5:0]    queue_3_exceptionInfo_eCode;
  reg        [0:0]    queue_3_exceptionInfo_eSubCode;
  reg        [31:0]   queue_3_pc;
  reg        [5:0]    queue_3_prd;
  reg        [5:0]    queue_3_psrc_0;
  reg        [5:0]    queue_3_psrc_1;
  reg        [31:0]   queue_3_imm;
  reg        [3:0]    queue_3_uop_lsuOp;
  reg        [4:0]    queue_3_uop_lsuCoOp;
  reg        [0:0]    queue_3_roop_lsuROOp;
  reg                 queue_3_srcReady_0;
  reg                 queue_3_srcReady_1;
  reg        [3:0]    readyToIssue;
  wire       [3:0]    readyToIssue_ohFirst_input;
  wire       [3:0]    readyToIssue_ohFirst_masked;
  wire       [3:0]    issueVector;
  reg        [3:0]    shiftAhead;
  reg        [4:0]    emptyEntry;
  wire       [4:0]    emptyEntry_ohFirst_input;
  wire       [4:0]    emptyEntry_ohFirst_masked;
  wire       [4:0]    writeVector;
  wire                updatedEntry_0_valid;
  wire       [4:0]    updatedEntry_0_robIdx;
  wire       [31:0]   updatedEntry_0_branchResult_targetPC;
  wire                updatedEntry_0_branchResult_branchResult;
  wire                updatedEntry_0_branchResult_predictFail;
  wire                updatedEntry_0_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_0_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_0_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_0_pc;
  wire       [5:0]    updatedEntry_0_prd;
  wire       [5:0]    updatedEntry_0_psrc_0;
  wire       [5:0]    updatedEntry_0_psrc_1;
  wire       [31:0]   updatedEntry_0_imm;
  wire       [3:0]    updatedEntry_0_uop_lsuOp;
  wire       [4:0]    updatedEntry_0_uop_lsuCoOp;
  wire       [0:0]    updatedEntry_0_roop_lsuROOp;
  reg                 updatedEntry_0_srcReady_0;
  reg                 updatedEntry_0_srcReady_1;
  wire                updatedEntry_1_valid;
  wire       [4:0]    updatedEntry_1_robIdx;
  wire       [31:0]   updatedEntry_1_branchResult_targetPC;
  wire                updatedEntry_1_branchResult_branchResult;
  wire                updatedEntry_1_branchResult_predictFail;
  wire                updatedEntry_1_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_1_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_1_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_1_pc;
  wire       [5:0]    updatedEntry_1_prd;
  wire       [5:0]    updatedEntry_1_psrc_0;
  wire       [5:0]    updatedEntry_1_psrc_1;
  wire       [31:0]   updatedEntry_1_imm;
  wire       [3:0]    updatedEntry_1_uop_lsuOp;
  wire       [4:0]    updatedEntry_1_uop_lsuCoOp;
  wire       [0:0]    updatedEntry_1_roop_lsuROOp;
  reg                 updatedEntry_1_srcReady_0;
  reg                 updatedEntry_1_srcReady_1;
  wire                updatedEntry_2_valid;
  wire       [4:0]    updatedEntry_2_robIdx;
  wire       [31:0]   updatedEntry_2_branchResult_targetPC;
  wire                updatedEntry_2_branchResult_branchResult;
  wire                updatedEntry_2_branchResult_predictFail;
  wire                updatedEntry_2_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_2_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_2_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_2_pc;
  wire       [5:0]    updatedEntry_2_prd;
  wire       [5:0]    updatedEntry_2_psrc_0;
  wire       [5:0]    updatedEntry_2_psrc_1;
  wire       [31:0]   updatedEntry_2_imm;
  wire       [3:0]    updatedEntry_2_uop_lsuOp;
  wire       [4:0]    updatedEntry_2_uop_lsuCoOp;
  wire       [0:0]    updatedEntry_2_roop_lsuROOp;
  reg                 updatedEntry_2_srcReady_0;
  reg                 updatedEntry_2_srcReady_1;
  wire                updatedEntry_3_valid;
  wire       [4:0]    updatedEntry_3_robIdx;
  wire       [31:0]   updatedEntry_3_branchResult_targetPC;
  wire                updatedEntry_3_branchResult_branchResult;
  wire                updatedEntry_3_branchResult_predictFail;
  wire                updatedEntry_3_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_3_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_3_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_3_pc;
  wire       [5:0]    updatedEntry_3_prd;
  wire       [5:0]    updatedEntry_3_psrc_0;
  wire       [5:0]    updatedEntry_3_psrc_1;
  wire       [31:0]   updatedEntry_3_imm;
  wire       [3:0]    updatedEntry_3_uop_lsuOp;
  wire       [4:0]    updatedEntry_3_uop_lsuCoOp;
  wire       [0:0]    updatedEntry_3_roop_lsuROOp;
  reg                 updatedEntry_3_srcReady_0;
  reg                 updatedEntry_3_srcReady_1;
  wire                appendEntry_valid;
  wire       [4:0]    appendEntry_robIdx;
  wire       [31:0]   appendEntry_branchResult_targetPC;
  wire                appendEntry_branchResult_branchResult;
  wire                appendEntry_branchResult_predictFail;
  wire                appendEntry_exceptionInfo_exception;
  wire       [5:0]    appendEntry_exceptionInfo_eCode;
  wire       [0:0]    appendEntry_exceptionInfo_eSubCode;
  wire       [31:0]   appendEntry_pc;
  wire       [5:0]    appendEntry_prd;
  wire       [5:0]    appendEntry_psrc_0;
  wire       [5:0]    appendEntry_psrc_1;
  wire       [31:0]   appendEntry_imm;
  wire       [3:0]    appendEntry_uop_lsuOp;
  wire       [4:0]    appendEntry_uop_lsuCoOp;
  wire       [0:0]    appendEntry_roop_lsuROOp;
  wire                appendEntry_srcReady_0;
  wire                appendEntry_srcReady_1;
  reg                 queueNext_0_valid;
  reg        [4:0]    queueNext_0_robIdx;
  reg        [31:0]   queueNext_0_branchResult_targetPC;
  reg                 queueNext_0_branchResult_branchResult;
  reg                 queueNext_0_branchResult_predictFail;
  reg                 queueNext_0_exceptionInfo_exception;
  reg        [5:0]    queueNext_0_exceptionInfo_eCode;
  reg        [0:0]    queueNext_0_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_0_pc;
  reg        [5:0]    queueNext_0_prd;
  reg        [5:0]    queueNext_0_psrc_0;
  reg        [5:0]    queueNext_0_psrc_1;
  reg        [31:0]   queueNext_0_imm;
  reg        [3:0]    queueNext_0_uop_lsuOp;
  reg        [4:0]    queueNext_0_uop_lsuCoOp;
  reg        [0:0]    queueNext_0_roop_lsuROOp;
  reg                 queueNext_0_srcReady_0;
  reg                 queueNext_0_srcReady_1;
  reg                 queueNext_1_valid;
  reg        [4:0]    queueNext_1_robIdx;
  reg        [31:0]   queueNext_1_branchResult_targetPC;
  reg                 queueNext_1_branchResult_branchResult;
  reg                 queueNext_1_branchResult_predictFail;
  reg                 queueNext_1_exceptionInfo_exception;
  reg        [5:0]    queueNext_1_exceptionInfo_eCode;
  reg        [0:0]    queueNext_1_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_1_pc;
  reg        [5:0]    queueNext_1_prd;
  reg        [5:0]    queueNext_1_psrc_0;
  reg        [5:0]    queueNext_1_psrc_1;
  reg        [31:0]   queueNext_1_imm;
  reg        [3:0]    queueNext_1_uop_lsuOp;
  reg        [4:0]    queueNext_1_uop_lsuCoOp;
  reg        [0:0]    queueNext_1_roop_lsuROOp;
  reg                 queueNext_1_srcReady_0;
  reg                 queueNext_1_srcReady_1;
  reg                 queueNext_2_valid;
  reg        [4:0]    queueNext_2_robIdx;
  reg        [31:0]   queueNext_2_branchResult_targetPC;
  reg                 queueNext_2_branchResult_branchResult;
  reg                 queueNext_2_branchResult_predictFail;
  reg                 queueNext_2_exceptionInfo_exception;
  reg        [5:0]    queueNext_2_exceptionInfo_eCode;
  reg        [0:0]    queueNext_2_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_2_pc;
  reg        [5:0]    queueNext_2_prd;
  reg        [5:0]    queueNext_2_psrc_0;
  reg        [5:0]    queueNext_2_psrc_1;
  reg        [31:0]   queueNext_2_imm;
  reg        [3:0]    queueNext_2_uop_lsuOp;
  reg        [4:0]    queueNext_2_uop_lsuCoOp;
  reg        [0:0]    queueNext_2_roop_lsuROOp;
  reg                 queueNext_2_srcReady_0;
  reg                 queueNext_2_srcReady_1;
  reg                 queueNext_3_valid;
  reg        [4:0]    queueNext_3_robIdx;
  reg        [31:0]   queueNext_3_branchResult_targetPC;
  reg                 queueNext_3_branchResult_branchResult;
  reg                 queueNext_3_branchResult_predictFail;
  reg                 queueNext_3_exceptionInfo_exception;
  reg        [5:0]    queueNext_3_exceptionInfo_eCode;
  reg        [0:0]    queueNext_3_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_3_pc;
  reg        [5:0]    queueNext_3_prd;
  reg        [5:0]    queueNext_3_psrc_0;
  reg        [5:0]    queueNext_3_psrc_1;
  reg        [31:0]   queueNext_3_imm;
  reg        [3:0]    queueNext_3_uop_lsuOp;
  reg        [4:0]    queueNext_3_uop_lsuCoOp;
  reg        [0:0]    queueNext_3_roop_lsuROOp;
  reg                 queueNext_3_srcReady_0;
  reg                 queueNext_3_srcReady_1;
  wire                when_IssueQueue_l81;
  wire                when_IssueQueue_l83;
  wire                when_IssueQueue_l96;
  wire                when_IssueQueue_l81_1;
  wire                when_IssueQueue_l83_1;
  wire                when_IssueQueue_l96_1;
  wire                when_IssueQueue_l81_2;
  wire                when_IssueQueue_l83_2;
  wire                when_IssueQueue_l96_2;
  wire                when_IssueQueue_l81_3;
  wire                when_IssueQueue_l89;
  wire                when_IssueQueue_l96_3;
  wire                io_output_fire;
  wire                _zz_issueEntry_valid;
  wire                _zz_issueEntry_valid_1;
  wire                _zz_issueEntry_valid_2;
  wire       [1:0]    _zz_issueEntry_valid_3;
  wire                issueEntry_valid;
  wire       [4:0]    issueEntry_robIdx;
  wire       [31:0]   issueEntry_branchResult_targetPC;
  wire                issueEntry_branchResult_branchResult;
  wire                issueEntry_branchResult_predictFail;
  wire                issueEntry_exceptionInfo_exception;
  wire       [5:0]    issueEntry_exceptionInfo_eCode;
  wire       [0:0]    issueEntry_exceptionInfo_eSubCode;
  wire       [31:0]   issueEntry_pc;
  wire       [5:0]    issueEntry_prd;
  wire       [5:0]    issueEntry_psrc_0;
  wire       [5:0]    issueEntry_psrc_1;
  wire       [31:0]   issueEntry_imm;
  wire       [3:0]    issueEntry_uop_lsuOp;
  wire       [4:0]    issueEntry_uop_lsuCoOp;
  wire       [0:0]    issueEntry_roop_lsuROOp;
  wire                issueEntry_srcReady_0;
  wire                issueEntry_srcReady_1;
  `ifndef SYNTHESIS
  reg [55:0] io_input_payload_uop_lsuOp_string;
  reg [47:0] io_input_payload_roop_lsuROOp_string;
  reg [55:0] io_output_payload_uop_lsuOp_string;
  reg [47:0] io_output_payload_roop_lsuROOp_string;
  reg [55:0] queue_0_uop_lsuOp_string;
  reg [47:0] queue_0_roop_lsuROOp_string;
  reg [55:0] queue_1_uop_lsuOp_string;
  reg [47:0] queue_1_roop_lsuROOp_string;
  reg [55:0] queue_2_uop_lsuOp_string;
  reg [47:0] queue_2_roop_lsuROOp_string;
  reg [55:0] queue_3_uop_lsuOp_string;
  reg [47:0] queue_3_roop_lsuROOp_string;
  reg [55:0] updatedEntry_0_uop_lsuOp_string;
  reg [47:0] updatedEntry_0_roop_lsuROOp_string;
  reg [55:0] updatedEntry_1_uop_lsuOp_string;
  reg [47:0] updatedEntry_1_roop_lsuROOp_string;
  reg [55:0] updatedEntry_2_uop_lsuOp_string;
  reg [47:0] updatedEntry_2_roop_lsuROOp_string;
  reg [55:0] updatedEntry_3_uop_lsuOp_string;
  reg [47:0] updatedEntry_3_roop_lsuROOp_string;
  reg [55:0] appendEntry_uop_lsuOp_string;
  reg [47:0] appendEntry_roop_lsuROOp_string;
  reg [55:0] queueNext_0_uop_lsuOp_string;
  reg [47:0] queueNext_0_roop_lsuROOp_string;
  reg [55:0] queueNext_1_uop_lsuOp_string;
  reg [47:0] queueNext_1_roop_lsuROOp_string;
  reg [55:0] queueNext_2_uop_lsuOp_string;
  reg [47:0] queueNext_2_roop_lsuROOp_string;
  reg [55:0] queueNext_3_uop_lsuOp_string;
  reg [47:0] queueNext_3_roop_lsuROOp_string;
  reg [55:0] issueEntry_uop_lsuOp_string;
  reg [47:0] issueEntry_roop_lsuROOp_string;
  `endif


  assign _zz_readyToIssue_ohFirst_masked = (readyToIssue_ohFirst_input - 4'b0001);
  assign _zz_emptyEntry_ohFirst_masked = (emptyEntry_ohFirst_input - 5'h01);
  assign _zz_appendEntry_srcReady_0 = (io_input_payload_psrc_0 == io_writebackSignal_3);
  assign _zz_appendEntry_srcReady_0_1 = (io_input_payload_psrc_0 == io_writebackSignal_2);
  assign _zz_appendEntry_srcReady_0_2 = {(io_input_payload_psrc_0 == io_writebackSignal_1),(io_input_payload_psrc_0 == io_writebackSignal_0)};
  assign _zz_appendEntry_srcReady_0_3 = (io_input_payload_psrc_0 == io_earlyWakeup_9_payload);
  assign _zz_appendEntry_srcReady_0_4 = ((io_input_payload_psrc_0 == io_earlyWakeup_8_payload) && io_earlyWakeup_8_valid);
  assign _zz_appendEntry_srcReady_0_5 = ((io_input_payload_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid);
  assign _zz_appendEntry_srcReady_0_6 = {((io_input_payload_psrc_0 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid),{(_zz_appendEntry_srcReady_0_7 && io_earlyWakeup_5_valid),{_zz_appendEntry_srcReady_0_8,{_zz_appendEntry_srcReady_0_9,_zz_appendEntry_srcReady_0_10}}}};
  assign _zz_appendEntry_srcReady_0_7 = (io_input_payload_psrc_0 == io_earlyWakeup_5_payload);
  assign _zz_appendEntry_srcReady_0_8 = ((io_input_payload_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_appendEntry_srcReady_0_9 = ((io_input_payload_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid);
  assign _zz_appendEntry_srcReady_0_10 = {((io_input_payload_psrc_0 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((io_input_payload_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((io_input_payload_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}};
  assign _zz_appendEntry_srcReady_1 = (io_input_payload_psrc_1 == io_writebackSignal_2);
  assign _zz_appendEntry_srcReady_1_1 = (io_input_payload_psrc_1 == io_writebackSignal_1);
  assign _zz_appendEntry_srcReady_1_2 = (io_input_payload_psrc_1 == io_writebackSignal_0);
  assign _zz_appendEntry_srcReady_1_3 = (io_input_payload_psrc_1 == io_earlyWakeup_8_payload);
  assign _zz_appendEntry_srcReady_1_4 = ((io_input_payload_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid);
  assign _zz_appendEntry_srcReady_1_5 = ((io_input_payload_psrc_1 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid);
  assign _zz_appendEntry_srcReady_1_6 = {((io_input_payload_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid),{((io_input_payload_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid),{(_zz_appendEntry_srcReady_1_7 && io_earlyWakeup_3_valid),{_zz_appendEntry_srcReady_1_8,{_zz_appendEntry_srcReady_1_9,_zz_appendEntry_srcReady_1_10}}}}};
  assign _zz_appendEntry_srcReady_1_7 = (io_input_payload_psrc_1 == io_earlyWakeup_3_payload);
  assign _zz_appendEntry_srcReady_1_8 = ((io_input_payload_psrc_1 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid);
  assign _zz_appendEntry_srcReady_1_9 = ((io_input_payload_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid);
  assign _zz_appendEntry_srcReady_1_10 = ((io_input_payload_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid);
  assign _zz_updatedEntry_0_srcReady_0 = (queue_0_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_0_srcReady_0_1 = (queue_0_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_0_srcReady_0_2 = (queue_0_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_0_srcReady_0_3 = (queue_0_psrc_0 == io_earlyWakeup_8_payload);
  assign _zz_updatedEntry_0_srcReady_0_4 = ((queue_0_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid);
  assign _zz_updatedEntry_0_srcReady_0_5 = ((queue_0_psrc_0 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid);
  assign _zz_updatedEntry_0_srcReady_0_6 = {((queue_0_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid),{((queue_0_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid),{((queue_0_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{(_zz_updatedEntry_0_srcReady_0_7 && io_earlyWakeup_2_valid),{_zz_updatedEntry_0_srcReady_0_8,_zz_updatedEntry_0_srcReady_0_9}}}}};
  assign _zz_updatedEntry_0_srcReady_0_7 = (queue_0_psrc_0 == io_earlyWakeup_2_payload);
  assign _zz_updatedEntry_0_srcReady_0_8 = ((queue_0_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid);
  assign _zz_updatedEntry_0_srcReady_0_9 = ((queue_0_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid);
  assign _zz_updatedEntry_0_srcReady_1 = (queue_0_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_0_srcReady_1_1 = (queue_0_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_0_srcReady_1_2 = (queue_0_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_0_srcReady_1_3 = (queue_0_psrc_1 == io_earlyWakeup_8_payload);
  assign _zz_updatedEntry_0_srcReady_1_4 = ((queue_0_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid);
  assign _zz_updatedEntry_0_srcReady_1_5 = ((queue_0_psrc_1 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid);
  assign _zz_updatedEntry_0_srcReady_1_6 = {((queue_0_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid),{((queue_0_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid),{((queue_0_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{(_zz_updatedEntry_0_srcReady_1_7 && io_earlyWakeup_2_valid),{_zz_updatedEntry_0_srcReady_1_8,_zz_updatedEntry_0_srcReady_1_9}}}}};
  assign _zz_updatedEntry_0_srcReady_1_7 = (queue_0_psrc_1 == io_earlyWakeup_2_payload);
  assign _zz_updatedEntry_0_srcReady_1_8 = ((queue_0_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid);
  assign _zz_updatedEntry_0_srcReady_1_9 = ((queue_0_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid);
  assign _zz_updatedEntry_1_srcReady_0 = (queue_1_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_1_srcReady_0_1 = (queue_1_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_1_srcReady_0_2 = (queue_1_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_1_srcReady_0_3 = (queue_1_psrc_0 == io_earlyWakeup_8_payload);
  assign _zz_updatedEntry_1_srcReady_0_4 = ((queue_1_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid);
  assign _zz_updatedEntry_1_srcReady_0_5 = ((queue_1_psrc_0 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid);
  assign _zz_updatedEntry_1_srcReady_0_6 = {((queue_1_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid),{((queue_1_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid),{((queue_1_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{(_zz_updatedEntry_1_srcReady_0_7 && io_earlyWakeup_2_valid),{_zz_updatedEntry_1_srcReady_0_8,_zz_updatedEntry_1_srcReady_0_9}}}}};
  assign _zz_updatedEntry_1_srcReady_0_7 = (queue_1_psrc_0 == io_earlyWakeup_2_payload);
  assign _zz_updatedEntry_1_srcReady_0_8 = ((queue_1_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid);
  assign _zz_updatedEntry_1_srcReady_0_9 = ((queue_1_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid);
  assign _zz_updatedEntry_1_srcReady_1 = (queue_1_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_1_srcReady_1_1 = (queue_1_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_1_srcReady_1_2 = (queue_1_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_1_srcReady_1_3 = (queue_1_psrc_1 == io_earlyWakeup_8_payload);
  assign _zz_updatedEntry_1_srcReady_1_4 = ((queue_1_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid);
  assign _zz_updatedEntry_1_srcReady_1_5 = ((queue_1_psrc_1 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid);
  assign _zz_updatedEntry_1_srcReady_1_6 = {((queue_1_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid),{((queue_1_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid),{((queue_1_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{(_zz_updatedEntry_1_srcReady_1_7 && io_earlyWakeup_2_valid),{_zz_updatedEntry_1_srcReady_1_8,_zz_updatedEntry_1_srcReady_1_9}}}}};
  assign _zz_updatedEntry_1_srcReady_1_7 = (queue_1_psrc_1 == io_earlyWakeup_2_payload);
  assign _zz_updatedEntry_1_srcReady_1_8 = ((queue_1_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid);
  assign _zz_updatedEntry_1_srcReady_1_9 = ((queue_1_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid);
  assign _zz_updatedEntry_2_srcReady_0 = (queue_2_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_2_srcReady_0_1 = (queue_2_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_2_srcReady_0_2 = (queue_2_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_2_srcReady_0_3 = (queue_2_psrc_0 == io_earlyWakeup_8_payload);
  assign _zz_updatedEntry_2_srcReady_0_4 = ((queue_2_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid);
  assign _zz_updatedEntry_2_srcReady_0_5 = ((queue_2_psrc_0 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid);
  assign _zz_updatedEntry_2_srcReady_0_6 = {((queue_2_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid),{((queue_2_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid),{((queue_2_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{(_zz_updatedEntry_2_srcReady_0_7 && io_earlyWakeup_2_valid),{_zz_updatedEntry_2_srcReady_0_8,_zz_updatedEntry_2_srcReady_0_9}}}}};
  assign _zz_updatedEntry_2_srcReady_0_7 = (queue_2_psrc_0 == io_earlyWakeup_2_payload);
  assign _zz_updatedEntry_2_srcReady_0_8 = ((queue_2_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid);
  assign _zz_updatedEntry_2_srcReady_0_9 = ((queue_2_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid);
  assign _zz_updatedEntry_2_srcReady_1 = (queue_2_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_2_srcReady_1_1 = (queue_2_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_2_srcReady_1_2 = (queue_2_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_2_srcReady_1_3 = (queue_2_psrc_1 == io_earlyWakeup_8_payload);
  assign _zz_updatedEntry_2_srcReady_1_4 = ((queue_2_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid);
  assign _zz_updatedEntry_2_srcReady_1_5 = ((queue_2_psrc_1 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid);
  assign _zz_updatedEntry_2_srcReady_1_6 = {((queue_2_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid),{((queue_2_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid),{((queue_2_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{(_zz_updatedEntry_2_srcReady_1_7 && io_earlyWakeup_2_valid),{_zz_updatedEntry_2_srcReady_1_8,_zz_updatedEntry_2_srcReady_1_9}}}}};
  assign _zz_updatedEntry_2_srcReady_1_7 = (queue_2_psrc_1 == io_earlyWakeup_2_payload);
  assign _zz_updatedEntry_2_srcReady_1_8 = ((queue_2_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid);
  assign _zz_updatedEntry_2_srcReady_1_9 = ((queue_2_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid);
  assign _zz_updatedEntry_3_srcReady_0 = (queue_3_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_3_srcReady_0_1 = (queue_3_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_3_srcReady_0_2 = (queue_3_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_3_srcReady_0_3 = (queue_3_psrc_0 == io_earlyWakeup_8_payload);
  assign _zz_updatedEntry_3_srcReady_0_4 = ((queue_3_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid);
  assign _zz_updatedEntry_3_srcReady_0_5 = ((queue_3_psrc_0 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid);
  assign _zz_updatedEntry_3_srcReady_0_6 = {((queue_3_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid),{((queue_3_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid),{((queue_3_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{(_zz_updatedEntry_3_srcReady_0_7 && io_earlyWakeup_2_valid),{_zz_updatedEntry_3_srcReady_0_8,_zz_updatedEntry_3_srcReady_0_9}}}}};
  assign _zz_updatedEntry_3_srcReady_0_7 = (queue_3_psrc_0 == io_earlyWakeup_2_payload);
  assign _zz_updatedEntry_3_srcReady_0_8 = ((queue_3_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid);
  assign _zz_updatedEntry_3_srcReady_0_9 = ((queue_3_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid);
  assign _zz_updatedEntry_3_srcReady_1 = (queue_3_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_3_srcReady_1_1 = (queue_3_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_3_srcReady_1_2 = (queue_3_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_3_srcReady_1_3 = (queue_3_psrc_1 == io_earlyWakeup_8_payload);
  assign _zz_updatedEntry_3_srcReady_1_4 = ((queue_3_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid);
  assign _zz_updatedEntry_3_srcReady_1_5 = ((queue_3_psrc_1 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid);
  assign _zz_updatedEntry_3_srcReady_1_6 = {((queue_3_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid),{((queue_3_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid),{((queue_3_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{(_zz_updatedEntry_3_srcReady_1_7 && io_earlyWakeup_2_valid),{_zz_updatedEntry_3_srcReady_1_8,_zz_updatedEntry_3_srcReady_1_9}}}}};
  assign _zz_updatedEntry_3_srcReady_1_7 = (queue_3_psrc_1 == io_earlyWakeup_2_payload);
  assign _zz_updatedEntry_3_srcReady_1_8 = ((queue_3_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid);
  assign _zz_updatedEntry_3_srcReady_1_9 = ((queue_3_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid);
  always @(*) begin
    case(_zz_issueEntry_valid_3)
      2'b00 : begin
        _zz_issueEntry_valid_4 = queue_0_valid;
        _zz_issueEntry_robIdx = queue_0_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_0_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_0_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_0_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_0_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_0_pc;
        _zz_issueEntry_prd = queue_0_prd;
        _zz_issueEntry_psrc_0 = queue_0_psrc_0;
        _zz_issueEntry_psrc_1 = queue_0_psrc_1;
        _zz_issueEntry_imm = queue_0_imm;
        _zz_issueEntry_uop_lsuOp = queue_0_uop_lsuOp;
        _zz_issueEntry_uop_lsuCoOp = queue_0_uop_lsuCoOp;
        _zz_issueEntry_roop_lsuROOp = queue_0_roop_lsuROOp;
        _zz_issueEntry_srcReady_0 = queue_0_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_0_srcReady_1;
      end
      2'b01 : begin
        _zz_issueEntry_valid_4 = queue_1_valid;
        _zz_issueEntry_robIdx = queue_1_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_1_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_1_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_1_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_1_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_1_pc;
        _zz_issueEntry_prd = queue_1_prd;
        _zz_issueEntry_psrc_0 = queue_1_psrc_0;
        _zz_issueEntry_psrc_1 = queue_1_psrc_1;
        _zz_issueEntry_imm = queue_1_imm;
        _zz_issueEntry_uop_lsuOp = queue_1_uop_lsuOp;
        _zz_issueEntry_uop_lsuCoOp = queue_1_uop_lsuCoOp;
        _zz_issueEntry_roop_lsuROOp = queue_1_roop_lsuROOp;
        _zz_issueEntry_srcReady_0 = queue_1_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_1_srcReady_1;
      end
      2'b10 : begin
        _zz_issueEntry_valid_4 = queue_2_valid;
        _zz_issueEntry_robIdx = queue_2_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_2_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_2_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_2_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_2_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_2_pc;
        _zz_issueEntry_prd = queue_2_prd;
        _zz_issueEntry_psrc_0 = queue_2_psrc_0;
        _zz_issueEntry_psrc_1 = queue_2_psrc_1;
        _zz_issueEntry_imm = queue_2_imm;
        _zz_issueEntry_uop_lsuOp = queue_2_uop_lsuOp;
        _zz_issueEntry_uop_lsuCoOp = queue_2_uop_lsuCoOp;
        _zz_issueEntry_roop_lsuROOp = queue_2_roop_lsuROOp;
        _zz_issueEntry_srcReady_0 = queue_2_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_2_srcReady_1;
      end
      default : begin
        _zz_issueEntry_valid_4 = queue_3_valid;
        _zz_issueEntry_robIdx = queue_3_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_3_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_3_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_3_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_3_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_3_pc;
        _zz_issueEntry_prd = queue_3_prd;
        _zz_issueEntry_psrc_0 = queue_3_psrc_0;
        _zz_issueEntry_psrc_1 = queue_3_psrc_1;
        _zz_issueEntry_imm = queue_3_imm;
        _zz_issueEntry_uop_lsuOp = queue_3_uop_lsuOp;
        _zz_issueEntry_uop_lsuCoOp = queue_3_uop_lsuCoOp;
        _zz_issueEntry_roop_lsuROOp = queue_3_roop_lsuROOp;
        _zz_issueEntry_srcReady_0 = queue_3_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_3_srcReady_1;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_uop_lsuOp)
      LSUOp_cacop : io_input_payload_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : io_input_payload_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : io_input_payload_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : io_input_payload_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : io_input_payload_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : io_input_payload_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : io_input_payload_uop_lsuOp_string = "ll     ";
      LSUOp_sc : io_input_payload_uop_lsuOp_string = "sc     ";
      LSUOp_ld : io_input_payload_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : io_input_payload_uop_lsuOp_string = "ldu    ";
      LSUOp_st : io_input_payload_uop_lsuOp_string = "st     ";
      LSUOp_preld : io_input_payload_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : io_input_payload_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : io_input_payload_uop_lsuOp_string = "ibar   ";
      default : io_input_payload_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_input_payload_roop_lsuROOp)
      LSUROOp_reg_1 : io_input_payload_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : io_input_payload_roop_lsuROOp_string = "regimm";
      default : io_input_payload_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_uop_lsuOp)
      LSUOp_cacop : io_output_payload_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : io_output_payload_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : io_output_payload_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : io_output_payload_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : io_output_payload_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : io_output_payload_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : io_output_payload_uop_lsuOp_string = "ll     ";
      LSUOp_sc : io_output_payload_uop_lsuOp_string = "sc     ";
      LSUOp_ld : io_output_payload_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : io_output_payload_uop_lsuOp_string = "ldu    ";
      LSUOp_st : io_output_payload_uop_lsuOp_string = "st     ";
      LSUOp_preld : io_output_payload_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : io_output_payload_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : io_output_payload_uop_lsuOp_string = "ibar   ";
      default : io_output_payload_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_roop_lsuROOp)
      LSUROOp_reg_1 : io_output_payload_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : io_output_payload_roop_lsuROOp_string = "regimm";
      default : io_output_payload_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queue_0_uop_lsuOp)
      LSUOp_cacop : queue_0_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : queue_0_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : queue_0_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : queue_0_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : queue_0_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : queue_0_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : queue_0_uop_lsuOp_string = "ll     ";
      LSUOp_sc : queue_0_uop_lsuOp_string = "sc     ";
      LSUOp_ld : queue_0_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : queue_0_uop_lsuOp_string = "ldu    ";
      LSUOp_st : queue_0_uop_lsuOp_string = "st     ";
      LSUOp_preld : queue_0_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : queue_0_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : queue_0_uop_lsuOp_string = "ibar   ";
      default : queue_0_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_0_roop_lsuROOp)
      LSUROOp_reg_1 : queue_0_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : queue_0_roop_lsuROOp_string = "regimm";
      default : queue_0_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queue_1_uop_lsuOp)
      LSUOp_cacop : queue_1_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : queue_1_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : queue_1_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : queue_1_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : queue_1_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : queue_1_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : queue_1_uop_lsuOp_string = "ll     ";
      LSUOp_sc : queue_1_uop_lsuOp_string = "sc     ";
      LSUOp_ld : queue_1_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : queue_1_uop_lsuOp_string = "ldu    ";
      LSUOp_st : queue_1_uop_lsuOp_string = "st     ";
      LSUOp_preld : queue_1_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : queue_1_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : queue_1_uop_lsuOp_string = "ibar   ";
      default : queue_1_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_1_roop_lsuROOp)
      LSUROOp_reg_1 : queue_1_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : queue_1_roop_lsuROOp_string = "regimm";
      default : queue_1_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queue_2_uop_lsuOp)
      LSUOp_cacop : queue_2_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : queue_2_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : queue_2_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : queue_2_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : queue_2_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : queue_2_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : queue_2_uop_lsuOp_string = "ll     ";
      LSUOp_sc : queue_2_uop_lsuOp_string = "sc     ";
      LSUOp_ld : queue_2_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : queue_2_uop_lsuOp_string = "ldu    ";
      LSUOp_st : queue_2_uop_lsuOp_string = "st     ";
      LSUOp_preld : queue_2_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : queue_2_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : queue_2_uop_lsuOp_string = "ibar   ";
      default : queue_2_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_2_roop_lsuROOp)
      LSUROOp_reg_1 : queue_2_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : queue_2_roop_lsuROOp_string = "regimm";
      default : queue_2_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queue_3_uop_lsuOp)
      LSUOp_cacop : queue_3_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : queue_3_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : queue_3_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : queue_3_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : queue_3_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : queue_3_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : queue_3_uop_lsuOp_string = "ll     ";
      LSUOp_sc : queue_3_uop_lsuOp_string = "sc     ";
      LSUOp_ld : queue_3_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : queue_3_uop_lsuOp_string = "ldu    ";
      LSUOp_st : queue_3_uop_lsuOp_string = "st     ";
      LSUOp_preld : queue_3_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : queue_3_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : queue_3_uop_lsuOp_string = "ibar   ";
      default : queue_3_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_3_roop_lsuROOp)
      LSUROOp_reg_1 : queue_3_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : queue_3_roop_lsuROOp_string = "regimm";
      default : queue_3_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_uop_lsuOp)
      LSUOp_cacop : updatedEntry_0_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : updatedEntry_0_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : updatedEntry_0_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : updatedEntry_0_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : updatedEntry_0_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : updatedEntry_0_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : updatedEntry_0_uop_lsuOp_string = "ll     ";
      LSUOp_sc : updatedEntry_0_uop_lsuOp_string = "sc     ";
      LSUOp_ld : updatedEntry_0_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : updatedEntry_0_uop_lsuOp_string = "ldu    ";
      LSUOp_st : updatedEntry_0_uop_lsuOp_string = "st     ";
      LSUOp_preld : updatedEntry_0_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : updatedEntry_0_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : updatedEntry_0_uop_lsuOp_string = "ibar   ";
      default : updatedEntry_0_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_roop_lsuROOp)
      LSUROOp_reg_1 : updatedEntry_0_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : updatedEntry_0_roop_lsuROOp_string = "regimm";
      default : updatedEntry_0_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_uop_lsuOp)
      LSUOp_cacop : updatedEntry_1_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : updatedEntry_1_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : updatedEntry_1_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : updatedEntry_1_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : updatedEntry_1_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : updatedEntry_1_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : updatedEntry_1_uop_lsuOp_string = "ll     ";
      LSUOp_sc : updatedEntry_1_uop_lsuOp_string = "sc     ";
      LSUOp_ld : updatedEntry_1_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : updatedEntry_1_uop_lsuOp_string = "ldu    ";
      LSUOp_st : updatedEntry_1_uop_lsuOp_string = "st     ";
      LSUOp_preld : updatedEntry_1_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : updatedEntry_1_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : updatedEntry_1_uop_lsuOp_string = "ibar   ";
      default : updatedEntry_1_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_roop_lsuROOp)
      LSUROOp_reg_1 : updatedEntry_1_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : updatedEntry_1_roop_lsuROOp_string = "regimm";
      default : updatedEntry_1_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_uop_lsuOp)
      LSUOp_cacop : updatedEntry_2_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : updatedEntry_2_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : updatedEntry_2_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : updatedEntry_2_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : updatedEntry_2_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : updatedEntry_2_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : updatedEntry_2_uop_lsuOp_string = "ll     ";
      LSUOp_sc : updatedEntry_2_uop_lsuOp_string = "sc     ";
      LSUOp_ld : updatedEntry_2_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : updatedEntry_2_uop_lsuOp_string = "ldu    ";
      LSUOp_st : updatedEntry_2_uop_lsuOp_string = "st     ";
      LSUOp_preld : updatedEntry_2_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : updatedEntry_2_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : updatedEntry_2_uop_lsuOp_string = "ibar   ";
      default : updatedEntry_2_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_roop_lsuROOp)
      LSUROOp_reg_1 : updatedEntry_2_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : updatedEntry_2_roop_lsuROOp_string = "regimm";
      default : updatedEntry_2_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_uop_lsuOp)
      LSUOp_cacop : updatedEntry_3_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : updatedEntry_3_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : updatedEntry_3_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : updatedEntry_3_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : updatedEntry_3_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : updatedEntry_3_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : updatedEntry_3_uop_lsuOp_string = "ll     ";
      LSUOp_sc : updatedEntry_3_uop_lsuOp_string = "sc     ";
      LSUOp_ld : updatedEntry_3_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : updatedEntry_3_uop_lsuOp_string = "ldu    ";
      LSUOp_st : updatedEntry_3_uop_lsuOp_string = "st     ";
      LSUOp_preld : updatedEntry_3_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : updatedEntry_3_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : updatedEntry_3_uop_lsuOp_string = "ibar   ";
      default : updatedEntry_3_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_roop_lsuROOp)
      LSUROOp_reg_1 : updatedEntry_3_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : updatedEntry_3_roop_lsuROOp_string = "regimm";
      default : updatedEntry_3_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(appendEntry_uop_lsuOp)
      LSUOp_cacop : appendEntry_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : appendEntry_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : appendEntry_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : appendEntry_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : appendEntry_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : appendEntry_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : appendEntry_uop_lsuOp_string = "ll     ";
      LSUOp_sc : appendEntry_uop_lsuOp_string = "sc     ";
      LSUOp_ld : appendEntry_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : appendEntry_uop_lsuOp_string = "ldu    ";
      LSUOp_st : appendEntry_uop_lsuOp_string = "st     ";
      LSUOp_preld : appendEntry_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : appendEntry_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : appendEntry_uop_lsuOp_string = "ibar   ";
      default : appendEntry_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(appendEntry_roop_lsuROOp)
      LSUROOp_reg_1 : appendEntry_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : appendEntry_roop_lsuROOp_string = "regimm";
      default : appendEntry_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queueNext_0_uop_lsuOp)
      LSUOp_cacop : queueNext_0_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : queueNext_0_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : queueNext_0_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : queueNext_0_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : queueNext_0_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : queueNext_0_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : queueNext_0_uop_lsuOp_string = "ll     ";
      LSUOp_sc : queueNext_0_uop_lsuOp_string = "sc     ";
      LSUOp_ld : queueNext_0_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : queueNext_0_uop_lsuOp_string = "ldu    ";
      LSUOp_st : queueNext_0_uop_lsuOp_string = "st     ";
      LSUOp_preld : queueNext_0_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : queueNext_0_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : queueNext_0_uop_lsuOp_string = "ibar   ";
      default : queueNext_0_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_0_roop_lsuROOp)
      LSUROOp_reg_1 : queueNext_0_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : queueNext_0_roop_lsuROOp_string = "regimm";
      default : queueNext_0_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queueNext_1_uop_lsuOp)
      LSUOp_cacop : queueNext_1_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : queueNext_1_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : queueNext_1_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : queueNext_1_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : queueNext_1_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : queueNext_1_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : queueNext_1_uop_lsuOp_string = "ll     ";
      LSUOp_sc : queueNext_1_uop_lsuOp_string = "sc     ";
      LSUOp_ld : queueNext_1_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : queueNext_1_uop_lsuOp_string = "ldu    ";
      LSUOp_st : queueNext_1_uop_lsuOp_string = "st     ";
      LSUOp_preld : queueNext_1_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : queueNext_1_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : queueNext_1_uop_lsuOp_string = "ibar   ";
      default : queueNext_1_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_1_roop_lsuROOp)
      LSUROOp_reg_1 : queueNext_1_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : queueNext_1_roop_lsuROOp_string = "regimm";
      default : queueNext_1_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queueNext_2_uop_lsuOp)
      LSUOp_cacop : queueNext_2_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : queueNext_2_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : queueNext_2_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : queueNext_2_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : queueNext_2_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : queueNext_2_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : queueNext_2_uop_lsuOp_string = "ll     ";
      LSUOp_sc : queueNext_2_uop_lsuOp_string = "sc     ";
      LSUOp_ld : queueNext_2_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : queueNext_2_uop_lsuOp_string = "ldu    ";
      LSUOp_st : queueNext_2_uop_lsuOp_string = "st     ";
      LSUOp_preld : queueNext_2_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : queueNext_2_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : queueNext_2_uop_lsuOp_string = "ibar   ";
      default : queueNext_2_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_2_roop_lsuROOp)
      LSUROOp_reg_1 : queueNext_2_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : queueNext_2_roop_lsuROOp_string = "regimm";
      default : queueNext_2_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queueNext_3_uop_lsuOp)
      LSUOp_cacop : queueNext_3_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : queueNext_3_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : queueNext_3_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : queueNext_3_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : queueNext_3_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : queueNext_3_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : queueNext_3_uop_lsuOp_string = "ll     ";
      LSUOp_sc : queueNext_3_uop_lsuOp_string = "sc     ";
      LSUOp_ld : queueNext_3_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : queueNext_3_uop_lsuOp_string = "ldu    ";
      LSUOp_st : queueNext_3_uop_lsuOp_string = "st     ";
      LSUOp_preld : queueNext_3_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : queueNext_3_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : queueNext_3_uop_lsuOp_string = "ibar   ";
      default : queueNext_3_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_3_roop_lsuROOp)
      LSUROOp_reg_1 : queueNext_3_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : queueNext_3_roop_lsuROOp_string = "regimm";
      default : queueNext_3_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(issueEntry_uop_lsuOp)
      LSUOp_cacop : issueEntry_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : issueEntry_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : issueEntry_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : issueEntry_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : issueEntry_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : issueEntry_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : issueEntry_uop_lsuOp_string = "ll     ";
      LSUOp_sc : issueEntry_uop_lsuOp_string = "sc     ";
      LSUOp_ld : issueEntry_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : issueEntry_uop_lsuOp_string = "ldu    ";
      LSUOp_st : issueEntry_uop_lsuOp_string = "st     ";
      LSUOp_preld : issueEntry_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : issueEntry_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : issueEntry_uop_lsuOp_string = "ibar   ";
      default : issueEntry_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(issueEntry_roop_lsuROOp)
      LSUROOp_reg_1 : issueEntry_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : issueEntry_roop_lsuROOp_string = "regimm";
      default : issueEntry_roop_lsuROOp_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    readyToIssue[0] = ((queue_0_valid && queue_0_srcReady_0) && queue_0_srcReady_1);
    readyToIssue[1] = 1'b0;
    readyToIssue[2] = 1'b0;
    readyToIssue[3] = 1'b0;
  end

  assign readyToIssue_ohFirst_input = readyToIssue;
  assign readyToIssue_ohFirst_masked = (readyToIssue_ohFirst_input & (~ _zz_readyToIssue_ohFirst_masked));
  assign issueVector = readyToIssue_ohFirst_masked;
  always @(*) begin
    emptyEntry[0] = (! queue_0_valid);
    emptyEntry[1] = (! queue_1_valid);
    emptyEntry[2] = (! queue_2_valid);
    emptyEntry[3] = (! queue_3_valid);
    emptyEntry[4] = 1'b1;
    emptyEntry[0] = (! queue_0_valid);
    emptyEntry[1] = (! queue_1_valid);
    emptyEntry[2] = (! queue_2_valid);
    emptyEntry[3] = (! queue_3_valid);
  end

  assign emptyEntry_ohFirst_input = emptyEntry;
  assign emptyEntry_ohFirst_masked = (emptyEntry_ohFirst_input & (~ _zz_emptyEntry_ohFirst_masked));
  assign writeVector = emptyEntry_ohFirst_masked;
  assign appendEntry_valid = io_input_valid;
  assign appendEntry_robIdx = io_input_payload_robIdx;
  assign appendEntry_branchResult_targetPC = io_input_payload_branchResult_targetPC;
  assign appendEntry_branchResult_branchResult = io_input_payload_branchResult_branchResult;
  assign appendEntry_branchResult_predictFail = io_input_payload_branchResult_predictFail;
  assign appendEntry_exceptionInfo_exception = io_input_payload_exceptionInfo_exception;
  assign appendEntry_exceptionInfo_eCode = io_input_payload_exceptionInfo_eCode;
  assign appendEntry_exceptionInfo_eSubCode = io_input_payload_exceptionInfo_eSubCode;
  assign appendEntry_pc = io_input_payload_pc;
  assign appendEntry_prd = io_input_payload_prd;
  assign appendEntry_psrc_0 = io_input_payload_psrc_0;
  assign appendEntry_psrc_1 = io_input_payload_psrc_1;
  assign appendEntry_imm = io_input_payload_imm;
  assign appendEntry_uop_lsuOp = io_input_payload_uop_lsuOp;
  assign appendEntry_uop_lsuCoOp = io_input_payload_uop_lsuCoOp;
  assign appendEntry_roop_lsuROOp = io_input_payload_roop_lsuROOp;
  assign appendEntry_srcReady_0 = ((io_input_payload_srcReady_0 || (|{(io_input_payload_psrc_0 == io_writebackSignal_4),{_zz_appendEntry_srcReady_0,{_zz_appendEntry_srcReady_0_1,_zz_appendEntry_srcReady_0_2}}})) || (|{((io_input_payload_psrc_0 == io_earlyWakeup_10_payload) && io_earlyWakeup_10_valid),{(_zz_appendEntry_srcReady_0_3 && io_earlyWakeup_9_valid),{_zz_appendEntry_srcReady_0_4,{_zz_appendEntry_srcReady_0_5,_zz_appendEntry_srcReady_0_6}}}}));
  assign appendEntry_srcReady_1 = ((io_input_payload_srcReady_1 || (|{(io_input_payload_psrc_1 == io_writebackSignal_4),{(io_input_payload_psrc_1 == io_writebackSignal_3),{_zz_appendEntry_srcReady_1,{_zz_appendEntry_srcReady_1_1,_zz_appendEntry_srcReady_1_2}}}})) || (|{((io_input_payload_psrc_1 == io_earlyWakeup_10_payload) && io_earlyWakeup_10_valid),{((io_input_payload_psrc_1 == io_earlyWakeup_9_payload) && io_earlyWakeup_9_valid),{(_zz_appendEntry_srcReady_1_3 && io_earlyWakeup_8_valid),{_zz_appendEntry_srcReady_1_4,{_zz_appendEntry_srcReady_1_5,_zz_appendEntry_srcReady_1_6}}}}}));
  assign updatedEntry_0_valid = queue_0_valid;
  assign updatedEntry_0_robIdx = queue_0_robIdx;
  assign updatedEntry_0_branchResult_targetPC = queue_0_branchResult_targetPC;
  assign updatedEntry_0_branchResult_branchResult = queue_0_branchResult_branchResult;
  assign updatedEntry_0_branchResult_predictFail = queue_0_branchResult_predictFail;
  assign updatedEntry_0_exceptionInfo_exception = queue_0_exceptionInfo_exception;
  assign updatedEntry_0_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
  assign updatedEntry_0_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
  assign updatedEntry_0_pc = queue_0_pc;
  assign updatedEntry_0_prd = queue_0_prd;
  assign updatedEntry_0_psrc_0 = queue_0_psrc_0;
  assign updatedEntry_0_psrc_1 = queue_0_psrc_1;
  assign updatedEntry_0_imm = queue_0_imm;
  assign updatedEntry_0_uop_lsuOp = queue_0_uop_lsuOp;
  assign updatedEntry_0_uop_lsuCoOp = queue_0_uop_lsuCoOp;
  assign updatedEntry_0_roop_lsuROOp = queue_0_roop_lsuROOp;
  always @(*) begin
    updatedEntry_0_srcReady_0 = queue_0_srcReady_0;
    updatedEntry_0_srcReady_0 = ((queue_0_srcReady_0 || (|{(queue_0_psrc_0 == io_writebackSignal_4),{(queue_0_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_0_srcReady_0,{_zz_updatedEntry_0_srcReady_0_1,_zz_updatedEntry_0_srcReady_0_2}}}})) || (|{((queue_0_psrc_0 == io_earlyWakeup_10_payload) && io_earlyWakeup_10_valid),{((queue_0_psrc_0 == io_earlyWakeup_9_payload) && io_earlyWakeup_9_valid),{(_zz_updatedEntry_0_srcReady_0_3 && io_earlyWakeup_8_valid),{_zz_updatedEntry_0_srcReady_0_4,{_zz_updatedEntry_0_srcReady_0_5,_zz_updatedEntry_0_srcReady_0_6}}}}}));
  end

  always @(*) begin
    updatedEntry_0_srcReady_1 = queue_0_srcReady_1;
    updatedEntry_0_srcReady_1 = ((queue_0_srcReady_1 || (|{(queue_0_psrc_1 == io_writebackSignal_4),{(queue_0_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_0_srcReady_1,{_zz_updatedEntry_0_srcReady_1_1,_zz_updatedEntry_0_srcReady_1_2}}}})) || (|{((queue_0_psrc_1 == io_earlyWakeup_10_payload) && io_earlyWakeup_10_valid),{((queue_0_psrc_1 == io_earlyWakeup_9_payload) && io_earlyWakeup_9_valid),{(_zz_updatedEntry_0_srcReady_1_3 && io_earlyWakeup_8_valid),{_zz_updatedEntry_0_srcReady_1_4,{_zz_updatedEntry_0_srcReady_1_5,_zz_updatedEntry_0_srcReady_1_6}}}}}));
  end

  assign updatedEntry_1_valid = queue_1_valid;
  assign updatedEntry_1_robIdx = queue_1_robIdx;
  assign updatedEntry_1_branchResult_targetPC = queue_1_branchResult_targetPC;
  assign updatedEntry_1_branchResult_branchResult = queue_1_branchResult_branchResult;
  assign updatedEntry_1_branchResult_predictFail = queue_1_branchResult_predictFail;
  assign updatedEntry_1_exceptionInfo_exception = queue_1_exceptionInfo_exception;
  assign updatedEntry_1_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
  assign updatedEntry_1_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
  assign updatedEntry_1_pc = queue_1_pc;
  assign updatedEntry_1_prd = queue_1_prd;
  assign updatedEntry_1_psrc_0 = queue_1_psrc_0;
  assign updatedEntry_1_psrc_1 = queue_1_psrc_1;
  assign updatedEntry_1_imm = queue_1_imm;
  assign updatedEntry_1_uop_lsuOp = queue_1_uop_lsuOp;
  assign updatedEntry_1_uop_lsuCoOp = queue_1_uop_lsuCoOp;
  assign updatedEntry_1_roop_lsuROOp = queue_1_roop_lsuROOp;
  always @(*) begin
    updatedEntry_1_srcReady_0 = queue_1_srcReady_0;
    updatedEntry_1_srcReady_0 = ((queue_1_srcReady_0 || (|{(queue_1_psrc_0 == io_writebackSignal_4),{(queue_1_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_1_srcReady_0,{_zz_updatedEntry_1_srcReady_0_1,_zz_updatedEntry_1_srcReady_0_2}}}})) || (|{((queue_1_psrc_0 == io_earlyWakeup_10_payload) && io_earlyWakeup_10_valid),{((queue_1_psrc_0 == io_earlyWakeup_9_payload) && io_earlyWakeup_9_valid),{(_zz_updatedEntry_1_srcReady_0_3 && io_earlyWakeup_8_valid),{_zz_updatedEntry_1_srcReady_0_4,{_zz_updatedEntry_1_srcReady_0_5,_zz_updatedEntry_1_srcReady_0_6}}}}}));
  end

  always @(*) begin
    updatedEntry_1_srcReady_1 = queue_1_srcReady_1;
    updatedEntry_1_srcReady_1 = ((queue_1_srcReady_1 || (|{(queue_1_psrc_1 == io_writebackSignal_4),{(queue_1_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_1_srcReady_1,{_zz_updatedEntry_1_srcReady_1_1,_zz_updatedEntry_1_srcReady_1_2}}}})) || (|{((queue_1_psrc_1 == io_earlyWakeup_10_payload) && io_earlyWakeup_10_valid),{((queue_1_psrc_1 == io_earlyWakeup_9_payload) && io_earlyWakeup_9_valid),{(_zz_updatedEntry_1_srcReady_1_3 && io_earlyWakeup_8_valid),{_zz_updatedEntry_1_srcReady_1_4,{_zz_updatedEntry_1_srcReady_1_5,_zz_updatedEntry_1_srcReady_1_6}}}}}));
  end

  assign updatedEntry_2_valid = queue_2_valid;
  assign updatedEntry_2_robIdx = queue_2_robIdx;
  assign updatedEntry_2_branchResult_targetPC = queue_2_branchResult_targetPC;
  assign updatedEntry_2_branchResult_branchResult = queue_2_branchResult_branchResult;
  assign updatedEntry_2_branchResult_predictFail = queue_2_branchResult_predictFail;
  assign updatedEntry_2_exceptionInfo_exception = queue_2_exceptionInfo_exception;
  assign updatedEntry_2_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
  assign updatedEntry_2_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
  assign updatedEntry_2_pc = queue_2_pc;
  assign updatedEntry_2_prd = queue_2_prd;
  assign updatedEntry_2_psrc_0 = queue_2_psrc_0;
  assign updatedEntry_2_psrc_1 = queue_2_psrc_1;
  assign updatedEntry_2_imm = queue_2_imm;
  assign updatedEntry_2_uop_lsuOp = queue_2_uop_lsuOp;
  assign updatedEntry_2_uop_lsuCoOp = queue_2_uop_lsuCoOp;
  assign updatedEntry_2_roop_lsuROOp = queue_2_roop_lsuROOp;
  always @(*) begin
    updatedEntry_2_srcReady_0 = queue_2_srcReady_0;
    updatedEntry_2_srcReady_0 = ((queue_2_srcReady_0 || (|{(queue_2_psrc_0 == io_writebackSignal_4),{(queue_2_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_2_srcReady_0,{_zz_updatedEntry_2_srcReady_0_1,_zz_updatedEntry_2_srcReady_0_2}}}})) || (|{((queue_2_psrc_0 == io_earlyWakeup_10_payload) && io_earlyWakeup_10_valid),{((queue_2_psrc_0 == io_earlyWakeup_9_payload) && io_earlyWakeup_9_valid),{(_zz_updatedEntry_2_srcReady_0_3 && io_earlyWakeup_8_valid),{_zz_updatedEntry_2_srcReady_0_4,{_zz_updatedEntry_2_srcReady_0_5,_zz_updatedEntry_2_srcReady_0_6}}}}}));
  end

  always @(*) begin
    updatedEntry_2_srcReady_1 = queue_2_srcReady_1;
    updatedEntry_2_srcReady_1 = ((queue_2_srcReady_1 || (|{(queue_2_psrc_1 == io_writebackSignal_4),{(queue_2_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_2_srcReady_1,{_zz_updatedEntry_2_srcReady_1_1,_zz_updatedEntry_2_srcReady_1_2}}}})) || (|{((queue_2_psrc_1 == io_earlyWakeup_10_payload) && io_earlyWakeup_10_valid),{((queue_2_psrc_1 == io_earlyWakeup_9_payload) && io_earlyWakeup_9_valid),{(_zz_updatedEntry_2_srcReady_1_3 && io_earlyWakeup_8_valid),{_zz_updatedEntry_2_srcReady_1_4,{_zz_updatedEntry_2_srcReady_1_5,_zz_updatedEntry_2_srcReady_1_6}}}}}));
  end

  assign updatedEntry_3_valid = queue_3_valid;
  assign updatedEntry_3_robIdx = queue_3_robIdx;
  assign updatedEntry_3_branchResult_targetPC = queue_3_branchResult_targetPC;
  assign updatedEntry_3_branchResult_branchResult = queue_3_branchResult_branchResult;
  assign updatedEntry_3_branchResult_predictFail = queue_3_branchResult_predictFail;
  assign updatedEntry_3_exceptionInfo_exception = queue_3_exceptionInfo_exception;
  assign updatedEntry_3_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
  assign updatedEntry_3_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
  assign updatedEntry_3_pc = queue_3_pc;
  assign updatedEntry_3_prd = queue_3_prd;
  assign updatedEntry_3_psrc_0 = queue_3_psrc_0;
  assign updatedEntry_3_psrc_1 = queue_3_psrc_1;
  assign updatedEntry_3_imm = queue_3_imm;
  assign updatedEntry_3_uop_lsuOp = queue_3_uop_lsuOp;
  assign updatedEntry_3_uop_lsuCoOp = queue_3_uop_lsuCoOp;
  assign updatedEntry_3_roop_lsuROOp = queue_3_roop_lsuROOp;
  always @(*) begin
    updatedEntry_3_srcReady_0 = queue_3_srcReady_0;
    updatedEntry_3_srcReady_0 = ((queue_3_srcReady_0 || (|{(queue_3_psrc_0 == io_writebackSignal_4),{(queue_3_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_3_srcReady_0,{_zz_updatedEntry_3_srcReady_0_1,_zz_updatedEntry_3_srcReady_0_2}}}})) || (|{((queue_3_psrc_0 == io_earlyWakeup_10_payload) && io_earlyWakeup_10_valid),{((queue_3_psrc_0 == io_earlyWakeup_9_payload) && io_earlyWakeup_9_valid),{(_zz_updatedEntry_3_srcReady_0_3 && io_earlyWakeup_8_valid),{_zz_updatedEntry_3_srcReady_0_4,{_zz_updatedEntry_3_srcReady_0_5,_zz_updatedEntry_3_srcReady_0_6}}}}}));
  end

  always @(*) begin
    updatedEntry_3_srcReady_1 = queue_3_srcReady_1;
    updatedEntry_3_srcReady_1 = ((queue_3_srcReady_1 || (|{(queue_3_psrc_1 == io_writebackSignal_4),{(queue_3_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_3_srcReady_1,{_zz_updatedEntry_3_srcReady_1_1,_zz_updatedEntry_3_srcReady_1_2}}}})) || (|{((queue_3_psrc_1 == io_earlyWakeup_10_payload) && io_earlyWakeup_10_valid),{((queue_3_psrc_1 == io_earlyWakeup_9_payload) && io_earlyWakeup_9_valid),{(_zz_updatedEntry_3_srcReady_1_3 && io_earlyWakeup_8_valid),{_zz_updatedEntry_3_srcReady_1_4,{_zz_updatedEntry_3_srcReady_1_5,_zz_updatedEntry_3_srcReady_1_6}}}}}));
  end

  always @(*) begin
    shiftAhead[0] = ((|readyToIssue[0 : 0]) && io_output_ready);
    shiftAhead[1] = ((|readyToIssue[1 : 0]) && io_output_ready);
    shiftAhead[2] = ((|readyToIssue[2 : 0]) && io_output_ready);
    shiftAhead[3] = ((|readyToIssue[3 : 0]) && io_output_ready);
  end

  assign when_IssueQueue_l81 = shiftAhead[0];
  assign when_IssueQueue_l83 = writeVector[1];
  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_valid = appendEntry_valid;
      end else begin
        queueNext_0_valid = queue_1_valid;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_valid = appendEntry_valid;
      end else begin
        queueNext_0_valid = queue_0_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_0_robIdx = queue_1_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_0_robIdx = queue_0_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_0_branchResult_targetPC = queue_1_branchResult_targetPC;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_0_branchResult_targetPC = queue_0_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_0_branchResult_branchResult = queue_1_branchResult_branchResult;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_0_branchResult_branchResult = queue_0_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_0_branchResult_predictFail = queue_1_branchResult_predictFail;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_0_branchResult_predictFail = queue_0_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_0_exceptionInfo_exception = queue_1_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_0_exceptionInfo_exception = queue_0_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_0_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_0_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_0_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_0_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_pc = appendEntry_pc;
      end else begin
        queueNext_0_pc = queue_1_pc;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_pc = appendEntry_pc;
      end else begin
        queueNext_0_pc = queue_0_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_prd = appendEntry_prd;
      end else begin
        queueNext_0_prd = queue_1_prd;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_prd = appendEntry_prd;
      end else begin
        queueNext_0_prd = queue_0_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_0_psrc_0 = queue_1_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_0_psrc_0 = queue_0_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_0_psrc_1 = queue_1_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_0_psrc_1 = queue_0_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_imm = appendEntry_imm;
      end else begin
        queueNext_0_imm = queue_1_imm;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_imm = appendEntry_imm;
      end else begin
        queueNext_0_imm = queue_0_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_uop_lsuOp = appendEntry_uop_lsuOp;
      end else begin
        queueNext_0_uop_lsuOp = queue_1_uop_lsuOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_uop_lsuOp = appendEntry_uop_lsuOp;
      end else begin
        queueNext_0_uop_lsuOp = queue_0_uop_lsuOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_uop_lsuCoOp = appendEntry_uop_lsuCoOp;
      end else begin
        queueNext_0_uop_lsuCoOp = queue_1_uop_lsuCoOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_uop_lsuCoOp = appendEntry_uop_lsuCoOp;
      end else begin
        queueNext_0_uop_lsuCoOp = queue_0_uop_lsuCoOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_roop_lsuROOp = appendEntry_roop_lsuROOp;
      end else begin
        queueNext_0_roop_lsuROOp = queue_1_roop_lsuROOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_roop_lsuROOp = appendEntry_roop_lsuROOp;
      end else begin
        queueNext_0_roop_lsuROOp = queue_0_roop_lsuROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_0_srcReady_0 = queue_1_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_0_srcReady_0 = queue_0_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_0_srcReady_1 = queue_1_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_0_srcReady_1 = queue_0_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96 = writeVector[0];
  assign when_IssueQueue_l81_1 = shiftAhead[1];
  assign when_IssueQueue_l83_1 = writeVector[2];
  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_valid = appendEntry_valid;
      end else begin
        queueNext_1_valid = queue_2_valid;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_valid = appendEntry_valid;
      end else begin
        queueNext_1_valid = queue_1_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_1_robIdx = queue_2_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_1_robIdx = queue_1_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_1_branchResult_targetPC = queue_2_branchResult_targetPC;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_1_branchResult_targetPC = queue_1_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_1_branchResult_branchResult = queue_2_branchResult_branchResult;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_1_branchResult_branchResult = queue_1_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_1_branchResult_predictFail = queue_2_branchResult_predictFail;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_1_branchResult_predictFail = queue_1_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_1_exceptionInfo_exception = queue_2_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_1_exceptionInfo_exception = queue_1_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_1_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_1_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_1_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_1_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_pc = appendEntry_pc;
      end else begin
        queueNext_1_pc = queue_2_pc;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_pc = appendEntry_pc;
      end else begin
        queueNext_1_pc = queue_1_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_prd = appendEntry_prd;
      end else begin
        queueNext_1_prd = queue_2_prd;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_prd = appendEntry_prd;
      end else begin
        queueNext_1_prd = queue_1_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_1_psrc_0 = queue_2_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_1_psrc_0 = queue_1_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_1_psrc_1 = queue_2_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_1_psrc_1 = queue_1_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_imm = appendEntry_imm;
      end else begin
        queueNext_1_imm = queue_2_imm;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_imm = appendEntry_imm;
      end else begin
        queueNext_1_imm = queue_1_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_uop_lsuOp = appendEntry_uop_lsuOp;
      end else begin
        queueNext_1_uop_lsuOp = queue_2_uop_lsuOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_uop_lsuOp = appendEntry_uop_lsuOp;
      end else begin
        queueNext_1_uop_lsuOp = queue_1_uop_lsuOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_uop_lsuCoOp = appendEntry_uop_lsuCoOp;
      end else begin
        queueNext_1_uop_lsuCoOp = queue_2_uop_lsuCoOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_uop_lsuCoOp = appendEntry_uop_lsuCoOp;
      end else begin
        queueNext_1_uop_lsuCoOp = queue_1_uop_lsuCoOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_roop_lsuROOp = appendEntry_roop_lsuROOp;
      end else begin
        queueNext_1_roop_lsuROOp = queue_2_roop_lsuROOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_roop_lsuROOp = appendEntry_roop_lsuROOp;
      end else begin
        queueNext_1_roop_lsuROOp = queue_1_roop_lsuROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_1_srcReady_0 = queue_2_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_1_srcReady_0 = queue_1_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_1_srcReady_1 = queue_2_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_1_srcReady_1 = queue_1_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_1 = writeVector[1];
  assign when_IssueQueue_l81_2 = shiftAhead[2];
  assign when_IssueQueue_l83_2 = writeVector[3];
  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_valid = appendEntry_valid;
      end else begin
        queueNext_2_valid = queue_3_valid;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_valid = appendEntry_valid;
      end else begin
        queueNext_2_valid = queue_2_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_2_robIdx = queue_3_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_2_robIdx = queue_2_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_2_branchResult_targetPC = queue_3_branchResult_targetPC;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_2_branchResult_targetPC = queue_2_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_2_branchResult_branchResult = queue_3_branchResult_branchResult;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_2_branchResult_branchResult = queue_2_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_2_branchResult_predictFail = queue_3_branchResult_predictFail;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_2_branchResult_predictFail = queue_2_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_2_exceptionInfo_exception = queue_3_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_2_exceptionInfo_exception = queue_2_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_2_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_2_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_2_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_2_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_pc = appendEntry_pc;
      end else begin
        queueNext_2_pc = queue_3_pc;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_pc = appendEntry_pc;
      end else begin
        queueNext_2_pc = queue_2_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_prd = appendEntry_prd;
      end else begin
        queueNext_2_prd = queue_3_prd;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_prd = appendEntry_prd;
      end else begin
        queueNext_2_prd = queue_2_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_2_psrc_0 = queue_3_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_2_psrc_0 = queue_2_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_2_psrc_1 = queue_3_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_2_psrc_1 = queue_2_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_imm = appendEntry_imm;
      end else begin
        queueNext_2_imm = queue_3_imm;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_imm = appendEntry_imm;
      end else begin
        queueNext_2_imm = queue_2_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_uop_lsuOp = appendEntry_uop_lsuOp;
      end else begin
        queueNext_2_uop_lsuOp = queue_3_uop_lsuOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_uop_lsuOp = appendEntry_uop_lsuOp;
      end else begin
        queueNext_2_uop_lsuOp = queue_2_uop_lsuOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_uop_lsuCoOp = appendEntry_uop_lsuCoOp;
      end else begin
        queueNext_2_uop_lsuCoOp = queue_3_uop_lsuCoOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_uop_lsuCoOp = appendEntry_uop_lsuCoOp;
      end else begin
        queueNext_2_uop_lsuCoOp = queue_2_uop_lsuCoOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_roop_lsuROOp = appendEntry_roop_lsuROOp;
      end else begin
        queueNext_2_roop_lsuROOp = queue_3_roop_lsuROOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_roop_lsuROOp = appendEntry_roop_lsuROOp;
      end else begin
        queueNext_2_roop_lsuROOp = queue_2_roop_lsuROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_2_srcReady_0 = queue_3_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_2_srcReady_0 = queue_2_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_2_srcReady_1 = queue_3_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_2_srcReady_1 = queue_2_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_2 = writeVector[2];
  assign when_IssueQueue_l81_3 = shiftAhead[3];
  assign when_IssueQueue_l89 = writeVector[4];
  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_valid = appendEntry_valid;
      end else begin
        queueNext_3_valid = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_valid = appendEntry_valid;
      end else begin
        queueNext_3_valid = queue_3_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_3_robIdx = 5'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_3_robIdx = queue_3_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_3_branchResult_targetPC = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_3_branchResult_targetPC = queue_3_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_3_branchResult_branchResult = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_3_branchResult_branchResult = queue_3_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_3_branchResult_predictFail = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_3_branchResult_predictFail = queue_3_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_3_exceptionInfo_exception = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_3_exceptionInfo_exception = queue_3_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_3_exceptionInfo_eCode = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_3_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_3_exceptionInfo_eSubCode = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_3_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_pc = appendEntry_pc;
      end else begin
        queueNext_3_pc = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_pc = appendEntry_pc;
      end else begin
        queueNext_3_pc = queue_3_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_prd = appendEntry_prd;
      end else begin
        queueNext_3_prd = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_prd = appendEntry_prd;
      end else begin
        queueNext_3_prd = queue_3_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_3_psrc_0 = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_3_psrc_0 = queue_3_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_3_psrc_1 = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_3_psrc_1 = queue_3_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_imm = appendEntry_imm;
      end else begin
        queueNext_3_imm = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_imm = appendEntry_imm;
      end else begin
        queueNext_3_imm = queue_3_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_uop_lsuOp = appendEntry_uop_lsuOp;
      end else begin
        queueNext_3_uop_lsuOp = LSUOp_dbar;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_uop_lsuOp = appendEntry_uop_lsuOp;
      end else begin
        queueNext_3_uop_lsuOp = queue_3_uop_lsuOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_uop_lsuCoOp = appendEntry_uop_lsuCoOp;
      end else begin
        queueNext_3_uop_lsuCoOp = 5'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_uop_lsuCoOp = appendEntry_uop_lsuCoOp;
      end else begin
        queueNext_3_uop_lsuCoOp = queue_3_uop_lsuCoOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_roop_lsuROOp = appendEntry_roop_lsuROOp;
      end else begin
        queueNext_3_roop_lsuROOp = LSUROOp_regimm;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_roop_lsuROOp = appendEntry_roop_lsuROOp;
      end else begin
        queueNext_3_roop_lsuROOp = queue_3_roop_lsuROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_3_srcReady_0 = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_3_srcReady_0 = queue_3_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_3_srcReady_1 = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_3_srcReady_1 = queue_3_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_3 = writeVector[3];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_input_ready = ((|emptyEntry[3 : 0]) || io_output_fire);
  assign _zz_issueEntry_valid = issueVector[3];
  assign _zz_issueEntry_valid_1 = (issueVector[1] || _zz_issueEntry_valid);
  assign _zz_issueEntry_valid_2 = (issueVector[2] || _zz_issueEntry_valid);
  assign _zz_issueEntry_valid_3 = {_zz_issueEntry_valid_2,_zz_issueEntry_valid_1};
  assign issueEntry_valid = _zz_issueEntry_valid_4;
  assign issueEntry_robIdx = _zz_issueEntry_robIdx;
  assign issueEntry_branchResult_targetPC = _zz_issueEntry_branchResult_targetPC;
  assign issueEntry_branchResult_branchResult = _zz_issueEntry_branchResult_branchResult;
  assign issueEntry_branchResult_predictFail = _zz_issueEntry_branchResult_predictFail;
  assign issueEntry_exceptionInfo_exception = _zz_issueEntry_exceptionInfo_exception;
  assign issueEntry_exceptionInfo_eCode = _zz_issueEntry_exceptionInfo_eCode;
  assign issueEntry_exceptionInfo_eSubCode = _zz_issueEntry_exceptionInfo_eSubCode;
  assign issueEntry_pc = _zz_issueEntry_pc;
  assign issueEntry_prd = _zz_issueEntry_prd;
  assign issueEntry_psrc_0 = _zz_issueEntry_psrc_0;
  assign issueEntry_psrc_1 = _zz_issueEntry_psrc_1;
  assign issueEntry_imm = _zz_issueEntry_imm;
  assign issueEntry_uop_lsuOp = _zz_issueEntry_uop_lsuOp;
  assign issueEntry_uop_lsuCoOp = _zz_issueEntry_uop_lsuCoOp;
  assign issueEntry_roop_lsuROOp = _zz_issueEntry_roop_lsuROOp;
  assign issueEntry_srcReady_0 = _zz_issueEntry_srcReady_0;
  assign issueEntry_srcReady_1 = _zz_issueEntry_srcReady_1;
  assign io_output_valid = (|readyToIssue);
  assign io_output_payload_robIdx = issueEntry_robIdx;
  assign io_output_payload_branchResult_targetPC = issueEntry_branchResult_targetPC;
  assign io_output_payload_branchResult_branchResult = issueEntry_branchResult_branchResult;
  assign io_output_payload_branchResult_predictFail = issueEntry_branchResult_predictFail;
  assign io_output_payload_exceptionInfo_exception = issueEntry_exceptionInfo_exception;
  assign io_output_payload_exceptionInfo_eCode = issueEntry_exceptionInfo_eCode;
  assign io_output_payload_exceptionInfo_eSubCode = issueEntry_exceptionInfo_eSubCode;
  assign io_output_payload_pc = issueEntry_pc;
  assign io_output_payload_prd = issueEntry_prd;
  assign io_output_payload_psrc_0 = issueEntry_psrc_0;
  assign io_output_payload_psrc_1 = issueEntry_psrc_1;
  assign io_output_payload_imm = issueEntry_imm;
  assign io_output_payload_uop_lsuOp = issueEntry_uop_lsuOp;
  assign io_output_payload_uop_lsuCoOp = issueEntry_uop_lsuCoOp;
  assign io_output_payload_roop_lsuROOp = issueEntry_roop_lsuROOp;
  always @(posedge aclk) begin
    if(!cpuClockingArea_areaFlushReset_newReset) begin
      queue_0_valid <= 1'b0;
      queue_0_robIdx <= 5'h00;
      queue_0_branchResult_targetPC <= 32'h00000000;
      queue_0_branchResult_branchResult <= 1'b0;
      queue_0_branchResult_predictFail <= 1'b0;
      queue_0_exceptionInfo_exception <= 1'b0;
      queue_0_exceptionInfo_eCode <= 6'h00;
      queue_0_exceptionInfo_eSubCode <= 1'b0;
      queue_0_pc <= 32'h00000000;
      queue_0_prd <= 6'h00;
      queue_0_psrc_0 <= 6'h00;
      queue_0_psrc_1 <= 6'h00;
      queue_0_imm <= 32'h00000000;
      queue_0_uop_lsuOp <= LSUOp_dbar;
      queue_0_uop_lsuCoOp <= 5'h00;
      queue_0_roop_lsuROOp <= LSUROOp_regimm;
      queue_0_srcReady_0 <= 1'b0;
      queue_0_srcReady_1 <= 1'b0;
      queue_1_valid <= 1'b0;
      queue_1_robIdx <= 5'h00;
      queue_1_branchResult_targetPC <= 32'h00000000;
      queue_1_branchResult_branchResult <= 1'b0;
      queue_1_branchResult_predictFail <= 1'b0;
      queue_1_exceptionInfo_exception <= 1'b0;
      queue_1_exceptionInfo_eCode <= 6'h00;
      queue_1_exceptionInfo_eSubCode <= 1'b0;
      queue_1_pc <= 32'h00000000;
      queue_1_prd <= 6'h00;
      queue_1_psrc_0 <= 6'h00;
      queue_1_psrc_1 <= 6'h00;
      queue_1_imm <= 32'h00000000;
      queue_1_uop_lsuOp <= LSUOp_dbar;
      queue_1_uop_lsuCoOp <= 5'h00;
      queue_1_roop_lsuROOp <= LSUROOp_regimm;
      queue_1_srcReady_0 <= 1'b0;
      queue_1_srcReady_1 <= 1'b0;
      queue_2_valid <= 1'b0;
      queue_2_robIdx <= 5'h00;
      queue_2_branchResult_targetPC <= 32'h00000000;
      queue_2_branchResult_branchResult <= 1'b0;
      queue_2_branchResult_predictFail <= 1'b0;
      queue_2_exceptionInfo_exception <= 1'b0;
      queue_2_exceptionInfo_eCode <= 6'h00;
      queue_2_exceptionInfo_eSubCode <= 1'b0;
      queue_2_pc <= 32'h00000000;
      queue_2_prd <= 6'h00;
      queue_2_psrc_0 <= 6'h00;
      queue_2_psrc_1 <= 6'h00;
      queue_2_imm <= 32'h00000000;
      queue_2_uop_lsuOp <= LSUOp_dbar;
      queue_2_uop_lsuCoOp <= 5'h00;
      queue_2_roop_lsuROOp <= LSUROOp_regimm;
      queue_2_srcReady_0 <= 1'b0;
      queue_2_srcReady_1 <= 1'b0;
      queue_3_valid <= 1'b0;
      queue_3_robIdx <= 5'h00;
      queue_3_branchResult_targetPC <= 32'h00000000;
      queue_3_branchResult_branchResult <= 1'b0;
      queue_3_branchResult_predictFail <= 1'b0;
      queue_3_exceptionInfo_exception <= 1'b0;
      queue_3_exceptionInfo_eCode <= 6'h00;
      queue_3_exceptionInfo_eSubCode <= 1'b0;
      queue_3_pc <= 32'h00000000;
      queue_3_prd <= 6'h00;
      queue_3_psrc_0 <= 6'h00;
      queue_3_psrc_1 <= 6'h00;
      queue_3_imm <= 32'h00000000;
      queue_3_uop_lsuOp <= LSUOp_dbar;
      queue_3_uop_lsuCoOp <= 5'h00;
      queue_3_roop_lsuROOp <= LSUROOp_regimm;
      queue_3_srcReady_0 <= 1'b0;
      queue_3_srcReady_1 <= 1'b0;
    end else begin
      queue_0_valid <= queueNext_0_valid;
      queue_0_robIdx <= queueNext_0_robIdx;
      queue_0_branchResult_targetPC <= queueNext_0_branchResult_targetPC;
      queue_0_branchResult_branchResult <= queueNext_0_branchResult_branchResult;
      queue_0_branchResult_predictFail <= queueNext_0_branchResult_predictFail;
      queue_0_exceptionInfo_exception <= queueNext_0_exceptionInfo_exception;
      queue_0_exceptionInfo_eCode <= queueNext_0_exceptionInfo_eCode;
      queue_0_exceptionInfo_eSubCode <= queueNext_0_exceptionInfo_eSubCode;
      queue_0_pc <= queueNext_0_pc;
      queue_0_prd <= queueNext_0_prd;
      queue_0_psrc_0 <= queueNext_0_psrc_0;
      queue_0_psrc_1 <= queueNext_0_psrc_1;
      queue_0_imm <= queueNext_0_imm;
      queue_0_uop_lsuOp <= queueNext_0_uop_lsuOp;
      queue_0_uop_lsuCoOp <= queueNext_0_uop_lsuCoOp;
      queue_0_roop_lsuROOp <= queueNext_0_roop_lsuROOp;
      queue_0_srcReady_0 <= queueNext_0_srcReady_0;
      queue_0_srcReady_1 <= queueNext_0_srcReady_1;
      queue_1_valid <= queueNext_1_valid;
      queue_1_robIdx <= queueNext_1_robIdx;
      queue_1_branchResult_targetPC <= queueNext_1_branchResult_targetPC;
      queue_1_branchResult_branchResult <= queueNext_1_branchResult_branchResult;
      queue_1_branchResult_predictFail <= queueNext_1_branchResult_predictFail;
      queue_1_exceptionInfo_exception <= queueNext_1_exceptionInfo_exception;
      queue_1_exceptionInfo_eCode <= queueNext_1_exceptionInfo_eCode;
      queue_1_exceptionInfo_eSubCode <= queueNext_1_exceptionInfo_eSubCode;
      queue_1_pc <= queueNext_1_pc;
      queue_1_prd <= queueNext_1_prd;
      queue_1_psrc_0 <= queueNext_1_psrc_0;
      queue_1_psrc_1 <= queueNext_1_psrc_1;
      queue_1_imm <= queueNext_1_imm;
      queue_1_uop_lsuOp <= queueNext_1_uop_lsuOp;
      queue_1_uop_lsuCoOp <= queueNext_1_uop_lsuCoOp;
      queue_1_roop_lsuROOp <= queueNext_1_roop_lsuROOp;
      queue_1_srcReady_0 <= queueNext_1_srcReady_0;
      queue_1_srcReady_1 <= queueNext_1_srcReady_1;
      queue_2_valid <= queueNext_2_valid;
      queue_2_robIdx <= queueNext_2_robIdx;
      queue_2_branchResult_targetPC <= queueNext_2_branchResult_targetPC;
      queue_2_branchResult_branchResult <= queueNext_2_branchResult_branchResult;
      queue_2_branchResult_predictFail <= queueNext_2_branchResult_predictFail;
      queue_2_exceptionInfo_exception <= queueNext_2_exceptionInfo_exception;
      queue_2_exceptionInfo_eCode <= queueNext_2_exceptionInfo_eCode;
      queue_2_exceptionInfo_eSubCode <= queueNext_2_exceptionInfo_eSubCode;
      queue_2_pc <= queueNext_2_pc;
      queue_2_prd <= queueNext_2_prd;
      queue_2_psrc_0 <= queueNext_2_psrc_0;
      queue_2_psrc_1 <= queueNext_2_psrc_1;
      queue_2_imm <= queueNext_2_imm;
      queue_2_uop_lsuOp <= queueNext_2_uop_lsuOp;
      queue_2_uop_lsuCoOp <= queueNext_2_uop_lsuCoOp;
      queue_2_roop_lsuROOp <= queueNext_2_roop_lsuROOp;
      queue_2_srcReady_0 <= queueNext_2_srcReady_0;
      queue_2_srcReady_1 <= queueNext_2_srcReady_1;
      queue_3_valid <= queueNext_3_valid;
      queue_3_robIdx <= queueNext_3_robIdx;
      queue_3_branchResult_targetPC <= queueNext_3_branchResult_targetPC;
      queue_3_branchResult_branchResult <= queueNext_3_branchResult_branchResult;
      queue_3_branchResult_predictFail <= queueNext_3_branchResult_predictFail;
      queue_3_exceptionInfo_exception <= queueNext_3_exceptionInfo_exception;
      queue_3_exceptionInfo_eCode <= queueNext_3_exceptionInfo_eCode;
      queue_3_exceptionInfo_eSubCode <= queueNext_3_exceptionInfo_eSubCode;
      queue_3_pc <= queueNext_3_pc;
      queue_3_prd <= queueNext_3_prd;
      queue_3_psrc_0 <= queueNext_3_psrc_0;
      queue_3_psrc_1 <= queueNext_3_psrc_1;
      queue_3_imm <= queueNext_3_imm;
      queue_3_uop_lsuOp <= queueNext_3_uop_lsuOp;
      queue_3_uop_lsuCoOp <= queueNext_3_uop_lsuCoOp;
      queue_3_roop_lsuROOp <= queueNext_3_roop_lsuROOp;
      queue_3_srcReady_0 <= queueNext_3_srcReady_0;
      queue_3_srcReady_1 <= queueNext_3_srcReady_1;
    end
  end


endmodule

module IssueQueue_3 (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [4:0]    io_input_payload_robIdx,
  input  wire [31:0]   io_input_payload_branchResult_targetPC,
  input  wire          io_input_payload_branchResult_branchResult,
  input  wire          io_input_payload_branchResult_predictFail,
  input  wire          io_input_payload_exceptionInfo_exception,
  input  wire [5:0]    io_input_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_input_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_payload_pc,
  input  wire [5:0]    io_input_payload_prd,
  input  wire [5:0]    io_input_payload_psrc_0,
  input  wire [5:0]    io_input_payload_psrc_1,
  input  wire [31:0]   io_input_payload_imm,
  input  wire [1:0]    io_input_payload_uop_divuOp,
  input  wire          io_input_payload_srcReady_0,
  input  wire          io_input_payload_srcReady_1,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [4:0]    io_output_payload_robIdx,
  output wire [31:0]   io_output_payload_branchResult_targetPC,
  output wire          io_output_payload_branchResult_branchResult,
  output wire          io_output_payload_branchResult_predictFail,
  output wire          io_output_payload_exceptionInfo_exception,
  output wire [5:0]    io_output_payload_exceptionInfo_eCode,
  output wire [0:0]    io_output_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_output_payload_pc,
  output wire [5:0]    io_output_payload_prd,
  output wire [5:0]    io_output_payload_psrc_0,
  output wire [5:0]    io_output_payload_psrc_1,
  output wire [31:0]   io_output_payload_imm,
  output wire [1:0]    io_output_payload_uop_divuOp,
  input  wire [5:0]    io_writebackSignal_0,
  input  wire [5:0]    io_writebackSignal_1,
  input  wire [5:0]    io_writebackSignal_2,
  input  wire [5:0]    io_writebackSignal_3,
  input  wire [5:0]    io_writebackSignal_4,
  input  wire          aclk,
  input  wire          cpuClockingArea_areaFlushReset_newReset
);
  localparam DIVUOp_div = 2'd0;
  localparam DIVUOp_divu = 2'd1;
  localparam DIVUOp_mod_1 = 2'd2;
  localparam DIVUOp_modu = 2'd3;

  wire       [3:0]    _zz_readyToIssue_ohFirst_masked;
  wire       [4:0]    _zz_emptyEntry_ohFirst_masked;
  reg                 _zz_issueEntry_valid_4;
  reg        [4:0]    _zz_issueEntry_robIdx;
  reg        [31:0]   _zz_issueEntry_branchResult_targetPC;
  reg                 _zz_issueEntry_branchResult_branchResult;
  reg                 _zz_issueEntry_branchResult_predictFail;
  reg                 _zz_issueEntry_exceptionInfo_exception;
  reg        [5:0]    _zz_issueEntry_exceptionInfo_eCode;
  reg        [0:0]    _zz_issueEntry_exceptionInfo_eSubCode;
  reg        [31:0]   _zz_issueEntry_pc;
  reg        [5:0]    _zz_issueEntry_prd;
  reg        [5:0]    _zz_issueEntry_psrc_0;
  reg        [5:0]    _zz_issueEntry_psrc_1;
  reg        [31:0]   _zz_issueEntry_imm;
  reg        [1:0]    _zz_issueEntry_uop_divuOp;
  reg                 _zz_issueEntry_srcReady_0;
  reg                 _zz_issueEntry_srcReady_1;
  reg                 queue_0_valid;
  reg        [4:0]    queue_0_robIdx;
  reg        [31:0]   queue_0_branchResult_targetPC;
  reg                 queue_0_branchResult_branchResult;
  reg                 queue_0_branchResult_predictFail;
  reg                 queue_0_exceptionInfo_exception;
  reg        [5:0]    queue_0_exceptionInfo_eCode;
  reg        [0:0]    queue_0_exceptionInfo_eSubCode;
  reg        [31:0]   queue_0_pc;
  reg        [5:0]    queue_0_prd;
  reg        [5:0]    queue_0_psrc_0;
  reg        [5:0]    queue_0_psrc_1;
  reg        [31:0]   queue_0_imm;
  reg        [1:0]    queue_0_uop_divuOp;
  reg                 queue_0_srcReady_0;
  reg                 queue_0_srcReady_1;
  reg                 queue_1_valid;
  reg        [4:0]    queue_1_robIdx;
  reg        [31:0]   queue_1_branchResult_targetPC;
  reg                 queue_1_branchResult_branchResult;
  reg                 queue_1_branchResult_predictFail;
  reg                 queue_1_exceptionInfo_exception;
  reg        [5:0]    queue_1_exceptionInfo_eCode;
  reg        [0:0]    queue_1_exceptionInfo_eSubCode;
  reg        [31:0]   queue_1_pc;
  reg        [5:0]    queue_1_prd;
  reg        [5:0]    queue_1_psrc_0;
  reg        [5:0]    queue_1_psrc_1;
  reg        [31:0]   queue_1_imm;
  reg        [1:0]    queue_1_uop_divuOp;
  reg                 queue_1_srcReady_0;
  reg                 queue_1_srcReady_1;
  reg                 queue_2_valid;
  reg        [4:0]    queue_2_robIdx;
  reg        [31:0]   queue_2_branchResult_targetPC;
  reg                 queue_2_branchResult_branchResult;
  reg                 queue_2_branchResult_predictFail;
  reg                 queue_2_exceptionInfo_exception;
  reg        [5:0]    queue_2_exceptionInfo_eCode;
  reg        [0:0]    queue_2_exceptionInfo_eSubCode;
  reg        [31:0]   queue_2_pc;
  reg        [5:0]    queue_2_prd;
  reg        [5:0]    queue_2_psrc_0;
  reg        [5:0]    queue_2_psrc_1;
  reg        [31:0]   queue_2_imm;
  reg        [1:0]    queue_2_uop_divuOp;
  reg                 queue_2_srcReady_0;
  reg                 queue_2_srcReady_1;
  reg                 queue_3_valid;
  reg        [4:0]    queue_3_robIdx;
  reg        [31:0]   queue_3_branchResult_targetPC;
  reg                 queue_3_branchResult_branchResult;
  reg                 queue_3_branchResult_predictFail;
  reg                 queue_3_exceptionInfo_exception;
  reg        [5:0]    queue_3_exceptionInfo_eCode;
  reg        [0:0]    queue_3_exceptionInfo_eSubCode;
  reg        [31:0]   queue_3_pc;
  reg        [5:0]    queue_3_prd;
  reg        [5:0]    queue_3_psrc_0;
  reg        [5:0]    queue_3_psrc_1;
  reg        [31:0]   queue_3_imm;
  reg        [1:0]    queue_3_uop_divuOp;
  reg                 queue_3_srcReady_0;
  reg                 queue_3_srcReady_1;
  reg        [3:0]    readyToIssue;
  wire       [3:0]    readyToIssue_ohFirst_input;
  wire       [3:0]    readyToIssue_ohFirst_masked;
  wire       [3:0]    issueVector;
  reg        [3:0]    shiftAhead;
  reg        [4:0]    emptyEntry;
  wire       [4:0]    emptyEntry_ohFirst_input;
  wire       [4:0]    emptyEntry_ohFirst_masked;
  wire       [4:0]    writeVector;
  wire                updatedEntry_0_valid;
  wire       [4:0]    updatedEntry_0_robIdx;
  wire       [31:0]   updatedEntry_0_branchResult_targetPC;
  wire                updatedEntry_0_branchResult_branchResult;
  wire                updatedEntry_0_branchResult_predictFail;
  wire                updatedEntry_0_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_0_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_0_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_0_pc;
  wire       [5:0]    updatedEntry_0_prd;
  wire       [5:0]    updatedEntry_0_psrc_0;
  wire       [5:0]    updatedEntry_0_psrc_1;
  wire       [31:0]   updatedEntry_0_imm;
  wire       [1:0]    updatedEntry_0_uop_divuOp;
  reg                 updatedEntry_0_srcReady_0;
  reg                 updatedEntry_0_srcReady_1;
  wire                updatedEntry_1_valid;
  wire       [4:0]    updatedEntry_1_robIdx;
  wire       [31:0]   updatedEntry_1_branchResult_targetPC;
  wire                updatedEntry_1_branchResult_branchResult;
  wire                updatedEntry_1_branchResult_predictFail;
  wire                updatedEntry_1_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_1_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_1_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_1_pc;
  wire       [5:0]    updatedEntry_1_prd;
  wire       [5:0]    updatedEntry_1_psrc_0;
  wire       [5:0]    updatedEntry_1_psrc_1;
  wire       [31:0]   updatedEntry_1_imm;
  wire       [1:0]    updatedEntry_1_uop_divuOp;
  reg                 updatedEntry_1_srcReady_0;
  reg                 updatedEntry_1_srcReady_1;
  wire                updatedEntry_2_valid;
  wire       [4:0]    updatedEntry_2_robIdx;
  wire       [31:0]   updatedEntry_2_branchResult_targetPC;
  wire                updatedEntry_2_branchResult_branchResult;
  wire                updatedEntry_2_branchResult_predictFail;
  wire                updatedEntry_2_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_2_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_2_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_2_pc;
  wire       [5:0]    updatedEntry_2_prd;
  wire       [5:0]    updatedEntry_2_psrc_0;
  wire       [5:0]    updatedEntry_2_psrc_1;
  wire       [31:0]   updatedEntry_2_imm;
  wire       [1:0]    updatedEntry_2_uop_divuOp;
  reg                 updatedEntry_2_srcReady_0;
  reg                 updatedEntry_2_srcReady_1;
  wire                updatedEntry_3_valid;
  wire       [4:0]    updatedEntry_3_robIdx;
  wire       [31:0]   updatedEntry_3_branchResult_targetPC;
  wire                updatedEntry_3_branchResult_branchResult;
  wire                updatedEntry_3_branchResult_predictFail;
  wire                updatedEntry_3_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_3_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_3_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_3_pc;
  wire       [5:0]    updatedEntry_3_prd;
  wire       [5:0]    updatedEntry_3_psrc_0;
  wire       [5:0]    updatedEntry_3_psrc_1;
  wire       [31:0]   updatedEntry_3_imm;
  wire       [1:0]    updatedEntry_3_uop_divuOp;
  reg                 updatedEntry_3_srcReady_0;
  reg                 updatedEntry_3_srcReady_1;
  wire                appendEntry_valid;
  wire       [4:0]    appendEntry_robIdx;
  wire       [31:0]   appendEntry_branchResult_targetPC;
  wire                appendEntry_branchResult_branchResult;
  wire                appendEntry_branchResult_predictFail;
  wire                appendEntry_exceptionInfo_exception;
  wire       [5:0]    appendEntry_exceptionInfo_eCode;
  wire       [0:0]    appendEntry_exceptionInfo_eSubCode;
  wire       [31:0]   appendEntry_pc;
  wire       [5:0]    appendEntry_prd;
  wire       [5:0]    appendEntry_psrc_0;
  wire       [5:0]    appendEntry_psrc_1;
  wire       [31:0]   appendEntry_imm;
  wire       [1:0]    appendEntry_uop_divuOp;
  wire                appendEntry_srcReady_0;
  wire                appendEntry_srcReady_1;
  reg                 queueNext_0_valid;
  reg        [4:0]    queueNext_0_robIdx;
  reg        [31:0]   queueNext_0_branchResult_targetPC;
  reg                 queueNext_0_branchResult_branchResult;
  reg                 queueNext_0_branchResult_predictFail;
  reg                 queueNext_0_exceptionInfo_exception;
  reg        [5:0]    queueNext_0_exceptionInfo_eCode;
  reg        [0:0]    queueNext_0_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_0_pc;
  reg        [5:0]    queueNext_0_prd;
  reg        [5:0]    queueNext_0_psrc_0;
  reg        [5:0]    queueNext_0_psrc_1;
  reg        [31:0]   queueNext_0_imm;
  reg        [1:0]    queueNext_0_uop_divuOp;
  reg                 queueNext_0_srcReady_0;
  reg                 queueNext_0_srcReady_1;
  reg                 queueNext_1_valid;
  reg        [4:0]    queueNext_1_robIdx;
  reg        [31:0]   queueNext_1_branchResult_targetPC;
  reg                 queueNext_1_branchResult_branchResult;
  reg                 queueNext_1_branchResult_predictFail;
  reg                 queueNext_1_exceptionInfo_exception;
  reg        [5:0]    queueNext_1_exceptionInfo_eCode;
  reg        [0:0]    queueNext_1_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_1_pc;
  reg        [5:0]    queueNext_1_prd;
  reg        [5:0]    queueNext_1_psrc_0;
  reg        [5:0]    queueNext_1_psrc_1;
  reg        [31:0]   queueNext_1_imm;
  reg        [1:0]    queueNext_1_uop_divuOp;
  reg                 queueNext_1_srcReady_0;
  reg                 queueNext_1_srcReady_1;
  reg                 queueNext_2_valid;
  reg        [4:0]    queueNext_2_robIdx;
  reg        [31:0]   queueNext_2_branchResult_targetPC;
  reg                 queueNext_2_branchResult_branchResult;
  reg                 queueNext_2_branchResult_predictFail;
  reg                 queueNext_2_exceptionInfo_exception;
  reg        [5:0]    queueNext_2_exceptionInfo_eCode;
  reg        [0:0]    queueNext_2_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_2_pc;
  reg        [5:0]    queueNext_2_prd;
  reg        [5:0]    queueNext_2_psrc_0;
  reg        [5:0]    queueNext_2_psrc_1;
  reg        [31:0]   queueNext_2_imm;
  reg        [1:0]    queueNext_2_uop_divuOp;
  reg                 queueNext_2_srcReady_0;
  reg                 queueNext_2_srcReady_1;
  reg                 queueNext_3_valid;
  reg        [4:0]    queueNext_3_robIdx;
  reg        [31:0]   queueNext_3_branchResult_targetPC;
  reg                 queueNext_3_branchResult_branchResult;
  reg                 queueNext_3_branchResult_predictFail;
  reg                 queueNext_3_exceptionInfo_exception;
  reg        [5:0]    queueNext_3_exceptionInfo_eCode;
  reg        [0:0]    queueNext_3_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_3_pc;
  reg        [5:0]    queueNext_3_prd;
  reg        [5:0]    queueNext_3_psrc_0;
  reg        [5:0]    queueNext_3_psrc_1;
  reg        [31:0]   queueNext_3_imm;
  reg        [1:0]    queueNext_3_uop_divuOp;
  reg                 queueNext_3_srcReady_0;
  reg                 queueNext_3_srcReady_1;
  wire                when_IssueQueue_l81;
  wire                when_IssueQueue_l83;
  wire                when_IssueQueue_l96;
  wire                when_IssueQueue_l81_1;
  wire                when_IssueQueue_l83_1;
  wire                when_IssueQueue_l96_1;
  wire                when_IssueQueue_l81_2;
  wire                when_IssueQueue_l83_2;
  wire                when_IssueQueue_l96_2;
  wire                when_IssueQueue_l81_3;
  wire                when_IssueQueue_l89;
  wire                when_IssueQueue_l96_3;
  wire                io_output_fire;
  wire                _zz_issueEntry_valid;
  wire                _zz_issueEntry_valid_1;
  wire                _zz_issueEntry_valid_2;
  wire       [1:0]    _zz_issueEntry_valid_3;
  wire                issueEntry_valid;
  wire       [4:0]    issueEntry_robIdx;
  wire       [31:0]   issueEntry_branchResult_targetPC;
  wire                issueEntry_branchResult_branchResult;
  wire                issueEntry_branchResult_predictFail;
  wire                issueEntry_exceptionInfo_exception;
  wire       [5:0]    issueEntry_exceptionInfo_eCode;
  wire       [0:0]    issueEntry_exceptionInfo_eSubCode;
  wire       [31:0]   issueEntry_pc;
  wire       [5:0]    issueEntry_prd;
  wire       [5:0]    issueEntry_psrc_0;
  wire       [5:0]    issueEntry_psrc_1;
  wire       [31:0]   issueEntry_imm;
  wire       [1:0]    issueEntry_uop_divuOp;
  wire                issueEntry_srcReady_0;
  wire                issueEntry_srcReady_1;
  `ifndef SYNTHESIS
  reg [39:0] io_input_payload_uop_divuOp_string;
  reg [39:0] io_output_payload_uop_divuOp_string;
  reg [39:0] queue_0_uop_divuOp_string;
  reg [39:0] queue_1_uop_divuOp_string;
  reg [39:0] queue_2_uop_divuOp_string;
  reg [39:0] queue_3_uop_divuOp_string;
  reg [39:0] updatedEntry_0_uop_divuOp_string;
  reg [39:0] updatedEntry_1_uop_divuOp_string;
  reg [39:0] updatedEntry_2_uop_divuOp_string;
  reg [39:0] updatedEntry_3_uop_divuOp_string;
  reg [39:0] appendEntry_uop_divuOp_string;
  reg [39:0] queueNext_0_uop_divuOp_string;
  reg [39:0] queueNext_1_uop_divuOp_string;
  reg [39:0] queueNext_2_uop_divuOp_string;
  reg [39:0] queueNext_3_uop_divuOp_string;
  reg [39:0] issueEntry_uop_divuOp_string;
  `endif


  assign _zz_readyToIssue_ohFirst_masked = (readyToIssue_ohFirst_input - 4'b0001);
  assign _zz_emptyEntry_ohFirst_masked = (emptyEntry_ohFirst_input - 5'h01);
  always @(*) begin
    case(_zz_issueEntry_valid_3)
      2'b00 : begin
        _zz_issueEntry_valid_4 = queue_0_valid;
        _zz_issueEntry_robIdx = queue_0_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_0_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_0_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_0_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_0_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_0_pc;
        _zz_issueEntry_prd = queue_0_prd;
        _zz_issueEntry_psrc_0 = queue_0_psrc_0;
        _zz_issueEntry_psrc_1 = queue_0_psrc_1;
        _zz_issueEntry_imm = queue_0_imm;
        _zz_issueEntry_uop_divuOp = queue_0_uop_divuOp;
        _zz_issueEntry_srcReady_0 = queue_0_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_0_srcReady_1;
      end
      2'b01 : begin
        _zz_issueEntry_valid_4 = queue_1_valid;
        _zz_issueEntry_robIdx = queue_1_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_1_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_1_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_1_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_1_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_1_pc;
        _zz_issueEntry_prd = queue_1_prd;
        _zz_issueEntry_psrc_0 = queue_1_psrc_0;
        _zz_issueEntry_psrc_1 = queue_1_psrc_1;
        _zz_issueEntry_imm = queue_1_imm;
        _zz_issueEntry_uop_divuOp = queue_1_uop_divuOp;
        _zz_issueEntry_srcReady_0 = queue_1_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_1_srcReady_1;
      end
      2'b10 : begin
        _zz_issueEntry_valid_4 = queue_2_valid;
        _zz_issueEntry_robIdx = queue_2_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_2_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_2_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_2_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_2_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_2_pc;
        _zz_issueEntry_prd = queue_2_prd;
        _zz_issueEntry_psrc_0 = queue_2_psrc_0;
        _zz_issueEntry_psrc_1 = queue_2_psrc_1;
        _zz_issueEntry_imm = queue_2_imm;
        _zz_issueEntry_uop_divuOp = queue_2_uop_divuOp;
        _zz_issueEntry_srcReady_0 = queue_2_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_2_srcReady_1;
      end
      default : begin
        _zz_issueEntry_valid_4 = queue_3_valid;
        _zz_issueEntry_robIdx = queue_3_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_3_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_3_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_3_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_3_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_3_pc;
        _zz_issueEntry_prd = queue_3_prd;
        _zz_issueEntry_psrc_0 = queue_3_psrc_0;
        _zz_issueEntry_psrc_1 = queue_3_psrc_1;
        _zz_issueEntry_imm = queue_3_imm;
        _zz_issueEntry_uop_divuOp = queue_3_uop_divuOp;
        _zz_issueEntry_srcReady_0 = queue_3_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_3_srcReady_1;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_uop_divuOp)
      DIVUOp_div : io_input_payload_uop_divuOp_string = "div  ";
      DIVUOp_divu : io_input_payload_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : io_input_payload_uop_divuOp_string = "mod_1";
      DIVUOp_modu : io_input_payload_uop_divuOp_string = "modu ";
      default : io_input_payload_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_uop_divuOp)
      DIVUOp_div : io_output_payload_uop_divuOp_string = "div  ";
      DIVUOp_divu : io_output_payload_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : io_output_payload_uop_divuOp_string = "mod_1";
      DIVUOp_modu : io_output_payload_uop_divuOp_string = "modu ";
      default : io_output_payload_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_0_uop_divuOp)
      DIVUOp_div : queue_0_uop_divuOp_string = "div  ";
      DIVUOp_divu : queue_0_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : queue_0_uop_divuOp_string = "mod_1";
      DIVUOp_modu : queue_0_uop_divuOp_string = "modu ";
      default : queue_0_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_1_uop_divuOp)
      DIVUOp_div : queue_1_uop_divuOp_string = "div  ";
      DIVUOp_divu : queue_1_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : queue_1_uop_divuOp_string = "mod_1";
      DIVUOp_modu : queue_1_uop_divuOp_string = "modu ";
      default : queue_1_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_2_uop_divuOp)
      DIVUOp_div : queue_2_uop_divuOp_string = "div  ";
      DIVUOp_divu : queue_2_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : queue_2_uop_divuOp_string = "mod_1";
      DIVUOp_modu : queue_2_uop_divuOp_string = "modu ";
      default : queue_2_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_3_uop_divuOp)
      DIVUOp_div : queue_3_uop_divuOp_string = "div  ";
      DIVUOp_divu : queue_3_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : queue_3_uop_divuOp_string = "mod_1";
      DIVUOp_modu : queue_3_uop_divuOp_string = "modu ";
      default : queue_3_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_uop_divuOp)
      DIVUOp_div : updatedEntry_0_uop_divuOp_string = "div  ";
      DIVUOp_divu : updatedEntry_0_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : updatedEntry_0_uop_divuOp_string = "mod_1";
      DIVUOp_modu : updatedEntry_0_uop_divuOp_string = "modu ";
      default : updatedEntry_0_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_uop_divuOp)
      DIVUOp_div : updatedEntry_1_uop_divuOp_string = "div  ";
      DIVUOp_divu : updatedEntry_1_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : updatedEntry_1_uop_divuOp_string = "mod_1";
      DIVUOp_modu : updatedEntry_1_uop_divuOp_string = "modu ";
      default : updatedEntry_1_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_uop_divuOp)
      DIVUOp_div : updatedEntry_2_uop_divuOp_string = "div  ";
      DIVUOp_divu : updatedEntry_2_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : updatedEntry_2_uop_divuOp_string = "mod_1";
      DIVUOp_modu : updatedEntry_2_uop_divuOp_string = "modu ";
      default : updatedEntry_2_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_uop_divuOp)
      DIVUOp_div : updatedEntry_3_uop_divuOp_string = "div  ";
      DIVUOp_divu : updatedEntry_3_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : updatedEntry_3_uop_divuOp_string = "mod_1";
      DIVUOp_modu : updatedEntry_3_uop_divuOp_string = "modu ";
      default : updatedEntry_3_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(appendEntry_uop_divuOp)
      DIVUOp_div : appendEntry_uop_divuOp_string = "div  ";
      DIVUOp_divu : appendEntry_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : appendEntry_uop_divuOp_string = "mod_1";
      DIVUOp_modu : appendEntry_uop_divuOp_string = "modu ";
      default : appendEntry_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_0_uop_divuOp)
      DIVUOp_div : queueNext_0_uop_divuOp_string = "div  ";
      DIVUOp_divu : queueNext_0_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : queueNext_0_uop_divuOp_string = "mod_1";
      DIVUOp_modu : queueNext_0_uop_divuOp_string = "modu ";
      default : queueNext_0_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_1_uop_divuOp)
      DIVUOp_div : queueNext_1_uop_divuOp_string = "div  ";
      DIVUOp_divu : queueNext_1_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : queueNext_1_uop_divuOp_string = "mod_1";
      DIVUOp_modu : queueNext_1_uop_divuOp_string = "modu ";
      default : queueNext_1_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_2_uop_divuOp)
      DIVUOp_div : queueNext_2_uop_divuOp_string = "div  ";
      DIVUOp_divu : queueNext_2_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : queueNext_2_uop_divuOp_string = "mod_1";
      DIVUOp_modu : queueNext_2_uop_divuOp_string = "modu ";
      default : queueNext_2_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_3_uop_divuOp)
      DIVUOp_div : queueNext_3_uop_divuOp_string = "div  ";
      DIVUOp_divu : queueNext_3_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : queueNext_3_uop_divuOp_string = "mod_1";
      DIVUOp_modu : queueNext_3_uop_divuOp_string = "modu ";
      default : queueNext_3_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(issueEntry_uop_divuOp)
      DIVUOp_div : issueEntry_uop_divuOp_string = "div  ";
      DIVUOp_divu : issueEntry_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : issueEntry_uop_divuOp_string = "mod_1";
      DIVUOp_modu : issueEntry_uop_divuOp_string = "modu ";
      default : issueEntry_uop_divuOp_string = "?????";
    endcase
  end
  `endif

  always @(*) begin
    readyToIssue[0] = (queue_0_valid && (&{queue_0_srcReady_1,queue_0_srcReady_0}));
    readyToIssue[1] = 1'b0;
    readyToIssue[2] = 1'b0;
    readyToIssue[3] = 1'b0;
  end

  assign readyToIssue_ohFirst_input = readyToIssue;
  assign readyToIssue_ohFirst_masked = (readyToIssue_ohFirst_input & (~ _zz_readyToIssue_ohFirst_masked));
  assign issueVector = readyToIssue_ohFirst_masked;
  always @(*) begin
    emptyEntry[0] = (! queue_0_valid);
    emptyEntry[1] = (! queue_1_valid);
    emptyEntry[2] = (! queue_2_valid);
    emptyEntry[3] = (! queue_3_valid);
    emptyEntry[4] = 1'b1;
    emptyEntry[0] = (! queue_0_valid);
    emptyEntry[1] = (! queue_1_valid);
    emptyEntry[2] = (! queue_2_valid);
    emptyEntry[3] = (! queue_3_valid);
  end

  assign emptyEntry_ohFirst_input = emptyEntry;
  assign emptyEntry_ohFirst_masked = (emptyEntry_ohFirst_input & (~ _zz_emptyEntry_ohFirst_masked));
  assign writeVector = emptyEntry_ohFirst_masked;
  assign appendEntry_valid = io_input_valid;
  assign appendEntry_robIdx = io_input_payload_robIdx;
  assign appendEntry_branchResult_targetPC = io_input_payload_branchResult_targetPC;
  assign appendEntry_branchResult_branchResult = io_input_payload_branchResult_branchResult;
  assign appendEntry_branchResult_predictFail = io_input_payload_branchResult_predictFail;
  assign appendEntry_exceptionInfo_exception = io_input_payload_exceptionInfo_exception;
  assign appendEntry_exceptionInfo_eCode = io_input_payload_exceptionInfo_eCode;
  assign appendEntry_exceptionInfo_eSubCode = io_input_payload_exceptionInfo_eSubCode;
  assign appendEntry_pc = io_input_payload_pc;
  assign appendEntry_prd = io_input_payload_prd;
  assign appendEntry_psrc_0 = io_input_payload_psrc_0;
  assign appendEntry_psrc_1 = io_input_payload_psrc_1;
  assign appendEntry_imm = io_input_payload_imm;
  assign appendEntry_uop_divuOp = io_input_payload_uop_divuOp;
  assign appendEntry_srcReady_0 = (io_input_payload_srcReady_0 || (|{(io_input_payload_psrc_0 == io_writebackSignal_4),{(io_input_payload_psrc_0 == io_writebackSignal_3),{(io_input_payload_psrc_0 == io_writebackSignal_2),{(io_input_payload_psrc_0 == io_writebackSignal_1),(io_input_payload_psrc_0 == io_writebackSignal_0)}}}}));
  assign appendEntry_srcReady_1 = (io_input_payload_srcReady_1 || (|{(io_input_payload_psrc_1 == io_writebackSignal_4),{(io_input_payload_psrc_1 == io_writebackSignal_3),{(io_input_payload_psrc_1 == io_writebackSignal_2),{(io_input_payload_psrc_1 == io_writebackSignal_1),(io_input_payload_psrc_1 == io_writebackSignal_0)}}}}));
  assign updatedEntry_0_valid = queue_0_valid;
  assign updatedEntry_0_robIdx = queue_0_robIdx;
  assign updatedEntry_0_branchResult_targetPC = queue_0_branchResult_targetPC;
  assign updatedEntry_0_branchResult_branchResult = queue_0_branchResult_branchResult;
  assign updatedEntry_0_branchResult_predictFail = queue_0_branchResult_predictFail;
  assign updatedEntry_0_exceptionInfo_exception = queue_0_exceptionInfo_exception;
  assign updatedEntry_0_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
  assign updatedEntry_0_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
  assign updatedEntry_0_pc = queue_0_pc;
  assign updatedEntry_0_prd = queue_0_prd;
  assign updatedEntry_0_psrc_0 = queue_0_psrc_0;
  assign updatedEntry_0_psrc_1 = queue_0_psrc_1;
  assign updatedEntry_0_imm = queue_0_imm;
  assign updatedEntry_0_uop_divuOp = queue_0_uop_divuOp;
  always @(*) begin
    updatedEntry_0_srcReady_0 = queue_0_srcReady_0;
    updatedEntry_0_srcReady_0 = (queue_0_srcReady_0 || (|{(queue_0_psrc_0 == io_writebackSignal_4),{(queue_0_psrc_0 == io_writebackSignal_3),{(queue_0_psrc_0 == io_writebackSignal_2),{(queue_0_psrc_0 == io_writebackSignal_1),(queue_0_psrc_0 == io_writebackSignal_0)}}}}));
  end

  always @(*) begin
    updatedEntry_0_srcReady_1 = queue_0_srcReady_1;
    updatedEntry_0_srcReady_1 = (queue_0_srcReady_1 || (|{(queue_0_psrc_1 == io_writebackSignal_4),{(queue_0_psrc_1 == io_writebackSignal_3),{(queue_0_psrc_1 == io_writebackSignal_2),{(queue_0_psrc_1 == io_writebackSignal_1),(queue_0_psrc_1 == io_writebackSignal_0)}}}}));
  end

  assign updatedEntry_1_valid = queue_1_valid;
  assign updatedEntry_1_robIdx = queue_1_robIdx;
  assign updatedEntry_1_branchResult_targetPC = queue_1_branchResult_targetPC;
  assign updatedEntry_1_branchResult_branchResult = queue_1_branchResult_branchResult;
  assign updatedEntry_1_branchResult_predictFail = queue_1_branchResult_predictFail;
  assign updatedEntry_1_exceptionInfo_exception = queue_1_exceptionInfo_exception;
  assign updatedEntry_1_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
  assign updatedEntry_1_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
  assign updatedEntry_1_pc = queue_1_pc;
  assign updatedEntry_1_prd = queue_1_prd;
  assign updatedEntry_1_psrc_0 = queue_1_psrc_0;
  assign updatedEntry_1_psrc_1 = queue_1_psrc_1;
  assign updatedEntry_1_imm = queue_1_imm;
  assign updatedEntry_1_uop_divuOp = queue_1_uop_divuOp;
  always @(*) begin
    updatedEntry_1_srcReady_0 = queue_1_srcReady_0;
    updatedEntry_1_srcReady_0 = (queue_1_srcReady_0 || (|{(queue_1_psrc_0 == io_writebackSignal_4),{(queue_1_psrc_0 == io_writebackSignal_3),{(queue_1_psrc_0 == io_writebackSignal_2),{(queue_1_psrc_0 == io_writebackSignal_1),(queue_1_psrc_0 == io_writebackSignal_0)}}}}));
  end

  always @(*) begin
    updatedEntry_1_srcReady_1 = queue_1_srcReady_1;
    updatedEntry_1_srcReady_1 = (queue_1_srcReady_1 || (|{(queue_1_psrc_1 == io_writebackSignal_4),{(queue_1_psrc_1 == io_writebackSignal_3),{(queue_1_psrc_1 == io_writebackSignal_2),{(queue_1_psrc_1 == io_writebackSignal_1),(queue_1_psrc_1 == io_writebackSignal_0)}}}}));
  end

  assign updatedEntry_2_valid = queue_2_valid;
  assign updatedEntry_2_robIdx = queue_2_robIdx;
  assign updatedEntry_2_branchResult_targetPC = queue_2_branchResult_targetPC;
  assign updatedEntry_2_branchResult_branchResult = queue_2_branchResult_branchResult;
  assign updatedEntry_2_branchResult_predictFail = queue_2_branchResult_predictFail;
  assign updatedEntry_2_exceptionInfo_exception = queue_2_exceptionInfo_exception;
  assign updatedEntry_2_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
  assign updatedEntry_2_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
  assign updatedEntry_2_pc = queue_2_pc;
  assign updatedEntry_2_prd = queue_2_prd;
  assign updatedEntry_2_psrc_0 = queue_2_psrc_0;
  assign updatedEntry_2_psrc_1 = queue_2_psrc_1;
  assign updatedEntry_2_imm = queue_2_imm;
  assign updatedEntry_2_uop_divuOp = queue_2_uop_divuOp;
  always @(*) begin
    updatedEntry_2_srcReady_0 = queue_2_srcReady_0;
    updatedEntry_2_srcReady_0 = (queue_2_srcReady_0 || (|{(queue_2_psrc_0 == io_writebackSignal_4),{(queue_2_psrc_0 == io_writebackSignal_3),{(queue_2_psrc_0 == io_writebackSignal_2),{(queue_2_psrc_0 == io_writebackSignal_1),(queue_2_psrc_0 == io_writebackSignal_0)}}}}));
  end

  always @(*) begin
    updatedEntry_2_srcReady_1 = queue_2_srcReady_1;
    updatedEntry_2_srcReady_1 = (queue_2_srcReady_1 || (|{(queue_2_psrc_1 == io_writebackSignal_4),{(queue_2_psrc_1 == io_writebackSignal_3),{(queue_2_psrc_1 == io_writebackSignal_2),{(queue_2_psrc_1 == io_writebackSignal_1),(queue_2_psrc_1 == io_writebackSignal_0)}}}}));
  end

  assign updatedEntry_3_valid = queue_3_valid;
  assign updatedEntry_3_robIdx = queue_3_robIdx;
  assign updatedEntry_3_branchResult_targetPC = queue_3_branchResult_targetPC;
  assign updatedEntry_3_branchResult_branchResult = queue_3_branchResult_branchResult;
  assign updatedEntry_3_branchResult_predictFail = queue_3_branchResult_predictFail;
  assign updatedEntry_3_exceptionInfo_exception = queue_3_exceptionInfo_exception;
  assign updatedEntry_3_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
  assign updatedEntry_3_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
  assign updatedEntry_3_pc = queue_3_pc;
  assign updatedEntry_3_prd = queue_3_prd;
  assign updatedEntry_3_psrc_0 = queue_3_psrc_0;
  assign updatedEntry_3_psrc_1 = queue_3_psrc_1;
  assign updatedEntry_3_imm = queue_3_imm;
  assign updatedEntry_3_uop_divuOp = queue_3_uop_divuOp;
  always @(*) begin
    updatedEntry_3_srcReady_0 = queue_3_srcReady_0;
    updatedEntry_3_srcReady_0 = (queue_3_srcReady_0 || (|{(queue_3_psrc_0 == io_writebackSignal_4),{(queue_3_psrc_0 == io_writebackSignal_3),{(queue_3_psrc_0 == io_writebackSignal_2),{(queue_3_psrc_0 == io_writebackSignal_1),(queue_3_psrc_0 == io_writebackSignal_0)}}}}));
  end

  always @(*) begin
    updatedEntry_3_srcReady_1 = queue_3_srcReady_1;
    updatedEntry_3_srcReady_1 = (queue_3_srcReady_1 || (|{(queue_3_psrc_1 == io_writebackSignal_4),{(queue_3_psrc_1 == io_writebackSignal_3),{(queue_3_psrc_1 == io_writebackSignal_2),{(queue_3_psrc_1 == io_writebackSignal_1),(queue_3_psrc_1 == io_writebackSignal_0)}}}}));
  end

  always @(*) begin
    shiftAhead[0] = ((|readyToIssue[0 : 0]) && io_output_ready);
    shiftAhead[1] = ((|readyToIssue[1 : 0]) && io_output_ready);
    shiftAhead[2] = ((|readyToIssue[2 : 0]) && io_output_ready);
    shiftAhead[3] = ((|readyToIssue[3 : 0]) && io_output_ready);
  end

  assign when_IssueQueue_l81 = shiftAhead[0];
  assign when_IssueQueue_l83 = writeVector[1];
  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_valid = appendEntry_valid;
      end else begin
        queueNext_0_valid = queue_1_valid;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_valid = appendEntry_valid;
      end else begin
        queueNext_0_valid = queue_0_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_0_robIdx = queue_1_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_0_robIdx = queue_0_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_0_branchResult_targetPC = queue_1_branchResult_targetPC;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_0_branchResult_targetPC = queue_0_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_0_branchResult_branchResult = queue_1_branchResult_branchResult;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_0_branchResult_branchResult = queue_0_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_0_branchResult_predictFail = queue_1_branchResult_predictFail;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_0_branchResult_predictFail = queue_0_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_0_exceptionInfo_exception = queue_1_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_0_exceptionInfo_exception = queue_0_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_0_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_0_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_0_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_0_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_pc = appendEntry_pc;
      end else begin
        queueNext_0_pc = queue_1_pc;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_pc = appendEntry_pc;
      end else begin
        queueNext_0_pc = queue_0_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_prd = appendEntry_prd;
      end else begin
        queueNext_0_prd = queue_1_prd;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_prd = appendEntry_prd;
      end else begin
        queueNext_0_prd = queue_0_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_0_psrc_0 = queue_1_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_0_psrc_0 = queue_0_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_0_psrc_1 = queue_1_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_0_psrc_1 = queue_0_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_imm = appendEntry_imm;
      end else begin
        queueNext_0_imm = queue_1_imm;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_imm = appendEntry_imm;
      end else begin
        queueNext_0_imm = queue_0_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_uop_divuOp = appendEntry_uop_divuOp;
      end else begin
        queueNext_0_uop_divuOp = queue_1_uop_divuOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_uop_divuOp = appendEntry_uop_divuOp;
      end else begin
        queueNext_0_uop_divuOp = queue_0_uop_divuOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_0_srcReady_0 = queue_1_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_0_srcReady_0 = queue_0_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_0_srcReady_1 = queue_1_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_0_srcReady_1 = queue_0_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96 = writeVector[0];
  assign when_IssueQueue_l81_1 = shiftAhead[1];
  assign when_IssueQueue_l83_1 = writeVector[2];
  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_valid = appendEntry_valid;
      end else begin
        queueNext_1_valid = queue_2_valid;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_valid = appendEntry_valid;
      end else begin
        queueNext_1_valid = queue_1_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_1_robIdx = queue_2_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_1_robIdx = queue_1_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_1_branchResult_targetPC = queue_2_branchResult_targetPC;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_1_branchResult_targetPC = queue_1_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_1_branchResult_branchResult = queue_2_branchResult_branchResult;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_1_branchResult_branchResult = queue_1_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_1_branchResult_predictFail = queue_2_branchResult_predictFail;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_1_branchResult_predictFail = queue_1_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_1_exceptionInfo_exception = queue_2_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_1_exceptionInfo_exception = queue_1_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_1_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_1_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_1_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_1_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_pc = appendEntry_pc;
      end else begin
        queueNext_1_pc = queue_2_pc;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_pc = appendEntry_pc;
      end else begin
        queueNext_1_pc = queue_1_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_prd = appendEntry_prd;
      end else begin
        queueNext_1_prd = queue_2_prd;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_prd = appendEntry_prd;
      end else begin
        queueNext_1_prd = queue_1_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_1_psrc_0 = queue_2_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_1_psrc_0 = queue_1_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_1_psrc_1 = queue_2_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_1_psrc_1 = queue_1_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_imm = appendEntry_imm;
      end else begin
        queueNext_1_imm = queue_2_imm;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_imm = appendEntry_imm;
      end else begin
        queueNext_1_imm = queue_1_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_uop_divuOp = appendEntry_uop_divuOp;
      end else begin
        queueNext_1_uop_divuOp = queue_2_uop_divuOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_uop_divuOp = appendEntry_uop_divuOp;
      end else begin
        queueNext_1_uop_divuOp = queue_1_uop_divuOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_1_srcReady_0 = queue_2_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_1_srcReady_0 = queue_1_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_1_srcReady_1 = queue_2_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_1_srcReady_1 = queue_1_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_1 = writeVector[1];
  assign when_IssueQueue_l81_2 = shiftAhead[2];
  assign when_IssueQueue_l83_2 = writeVector[3];
  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_valid = appendEntry_valid;
      end else begin
        queueNext_2_valid = queue_3_valid;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_valid = appendEntry_valid;
      end else begin
        queueNext_2_valid = queue_2_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_2_robIdx = queue_3_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_2_robIdx = queue_2_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_2_branchResult_targetPC = queue_3_branchResult_targetPC;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_2_branchResult_targetPC = queue_2_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_2_branchResult_branchResult = queue_3_branchResult_branchResult;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_2_branchResult_branchResult = queue_2_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_2_branchResult_predictFail = queue_3_branchResult_predictFail;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_2_branchResult_predictFail = queue_2_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_2_exceptionInfo_exception = queue_3_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_2_exceptionInfo_exception = queue_2_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_2_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_2_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_2_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_2_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_pc = appendEntry_pc;
      end else begin
        queueNext_2_pc = queue_3_pc;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_pc = appendEntry_pc;
      end else begin
        queueNext_2_pc = queue_2_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_prd = appendEntry_prd;
      end else begin
        queueNext_2_prd = queue_3_prd;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_prd = appendEntry_prd;
      end else begin
        queueNext_2_prd = queue_2_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_2_psrc_0 = queue_3_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_2_psrc_0 = queue_2_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_2_psrc_1 = queue_3_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_2_psrc_1 = queue_2_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_imm = appendEntry_imm;
      end else begin
        queueNext_2_imm = queue_3_imm;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_imm = appendEntry_imm;
      end else begin
        queueNext_2_imm = queue_2_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_uop_divuOp = appendEntry_uop_divuOp;
      end else begin
        queueNext_2_uop_divuOp = queue_3_uop_divuOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_uop_divuOp = appendEntry_uop_divuOp;
      end else begin
        queueNext_2_uop_divuOp = queue_2_uop_divuOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_2_srcReady_0 = queue_3_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_2_srcReady_0 = queue_2_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_2_srcReady_1 = queue_3_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_2_srcReady_1 = queue_2_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_2 = writeVector[2];
  assign when_IssueQueue_l81_3 = shiftAhead[3];
  assign when_IssueQueue_l89 = writeVector[4];
  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_valid = appendEntry_valid;
      end else begin
        queueNext_3_valid = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_valid = appendEntry_valid;
      end else begin
        queueNext_3_valid = queue_3_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_3_robIdx = 5'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_3_robIdx = queue_3_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_3_branchResult_targetPC = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_3_branchResult_targetPC = queue_3_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_3_branchResult_branchResult = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_3_branchResult_branchResult = queue_3_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_3_branchResult_predictFail = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_3_branchResult_predictFail = queue_3_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_3_exceptionInfo_exception = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_3_exceptionInfo_exception = queue_3_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_3_exceptionInfo_eCode = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_3_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_3_exceptionInfo_eSubCode = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_3_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_pc = appendEntry_pc;
      end else begin
        queueNext_3_pc = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_pc = appendEntry_pc;
      end else begin
        queueNext_3_pc = queue_3_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_prd = appendEntry_prd;
      end else begin
        queueNext_3_prd = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_prd = appendEntry_prd;
      end else begin
        queueNext_3_prd = queue_3_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_3_psrc_0 = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_3_psrc_0 = queue_3_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_3_psrc_1 = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_3_psrc_1 = queue_3_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_imm = appendEntry_imm;
      end else begin
        queueNext_3_imm = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_imm = appendEntry_imm;
      end else begin
        queueNext_3_imm = queue_3_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_uop_divuOp = appendEntry_uop_divuOp;
      end else begin
        queueNext_3_uop_divuOp = DIVUOp_div;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_uop_divuOp = appendEntry_uop_divuOp;
      end else begin
        queueNext_3_uop_divuOp = queue_3_uop_divuOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_3_srcReady_0 = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_3_srcReady_0 = queue_3_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_3_srcReady_1 = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_3_srcReady_1 = queue_3_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_3 = writeVector[3];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_input_ready = ((|emptyEntry[3 : 0]) || io_output_fire);
  assign _zz_issueEntry_valid = issueVector[3];
  assign _zz_issueEntry_valid_1 = (issueVector[1] || _zz_issueEntry_valid);
  assign _zz_issueEntry_valid_2 = (issueVector[2] || _zz_issueEntry_valid);
  assign _zz_issueEntry_valid_3 = {_zz_issueEntry_valid_2,_zz_issueEntry_valid_1};
  assign issueEntry_valid = _zz_issueEntry_valid_4;
  assign issueEntry_robIdx = _zz_issueEntry_robIdx;
  assign issueEntry_branchResult_targetPC = _zz_issueEntry_branchResult_targetPC;
  assign issueEntry_branchResult_branchResult = _zz_issueEntry_branchResult_branchResult;
  assign issueEntry_branchResult_predictFail = _zz_issueEntry_branchResult_predictFail;
  assign issueEntry_exceptionInfo_exception = _zz_issueEntry_exceptionInfo_exception;
  assign issueEntry_exceptionInfo_eCode = _zz_issueEntry_exceptionInfo_eCode;
  assign issueEntry_exceptionInfo_eSubCode = _zz_issueEntry_exceptionInfo_eSubCode;
  assign issueEntry_pc = _zz_issueEntry_pc;
  assign issueEntry_prd = _zz_issueEntry_prd;
  assign issueEntry_psrc_0 = _zz_issueEntry_psrc_0;
  assign issueEntry_psrc_1 = _zz_issueEntry_psrc_1;
  assign issueEntry_imm = _zz_issueEntry_imm;
  assign issueEntry_uop_divuOp = _zz_issueEntry_uop_divuOp;
  assign issueEntry_srcReady_0 = _zz_issueEntry_srcReady_0;
  assign issueEntry_srcReady_1 = _zz_issueEntry_srcReady_1;
  assign io_output_valid = (|readyToIssue);
  assign io_output_payload_robIdx = issueEntry_robIdx;
  assign io_output_payload_branchResult_targetPC = issueEntry_branchResult_targetPC;
  assign io_output_payload_branchResult_branchResult = issueEntry_branchResult_branchResult;
  assign io_output_payload_branchResult_predictFail = issueEntry_branchResult_predictFail;
  assign io_output_payload_exceptionInfo_exception = issueEntry_exceptionInfo_exception;
  assign io_output_payload_exceptionInfo_eCode = issueEntry_exceptionInfo_eCode;
  assign io_output_payload_exceptionInfo_eSubCode = issueEntry_exceptionInfo_eSubCode;
  assign io_output_payload_pc = issueEntry_pc;
  assign io_output_payload_prd = issueEntry_prd;
  assign io_output_payload_psrc_0 = issueEntry_psrc_0;
  assign io_output_payload_psrc_1 = issueEntry_psrc_1;
  assign io_output_payload_imm = issueEntry_imm;
  assign io_output_payload_uop_divuOp = issueEntry_uop_divuOp;
  always @(posedge aclk) begin
    if(!cpuClockingArea_areaFlushReset_newReset) begin
      queue_0_valid <= 1'b0;
      queue_0_robIdx <= 5'h00;
      queue_0_branchResult_targetPC <= 32'h00000000;
      queue_0_branchResult_branchResult <= 1'b0;
      queue_0_branchResult_predictFail <= 1'b0;
      queue_0_exceptionInfo_exception <= 1'b0;
      queue_0_exceptionInfo_eCode <= 6'h00;
      queue_0_exceptionInfo_eSubCode <= 1'b0;
      queue_0_pc <= 32'h00000000;
      queue_0_prd <= 6'h00;
      queue_0_psrc_0 <= 6'h00;
      queue_0_psrc_1 <= 6'h00;
      queue_0_imm <= 32'h00000000;
      queue_0_uop_divuOp <= DIVUOp_div;
      queue_0_srcReady_0 <= 1'b0;
      queue_0_srcReady_1 <= 1'b0;
      queue_1_valid <= 1'b0;
      queue_1_robIdx <= 5'h00;
      queue_1_branchResult_targetPC <= 32'h00000000;
      queue_1_branchResult_branchResult <= 1'b0;
      queue_1_branchResult_predictFail <= 1'b0;
      queue_1_exceptionInfo_exception <= 1'b0;
      queue_1_exceptionInfo_eCode <= 6'h00;
      queue_1_exceptionInfo_eSubCode <= 1'b0;
      queue_1_pc <= 32'h00000000;
      queue_1_prd <= 6'h00;
      queue_1_psrc_0 <= 6'h00;
      queue_1_psrc_1 <= 6'h00;
      queue_1_imm <= 32'h00000000;
      queue_1_uop_divuOp <= DIVUOp_div;
      queue_1_srcReady_0 <= 1'b0;
      queue_1_srcReady_1 <= 1'b0;
      queue_2_valid <= 1'b0;
      queue_2_robIdx <= 5'h00;
      queue_2_branchResult_targetPC <= 32'h00000000;
      queue_2_branchResult_branchResult <= 1'b0;
      queue_2_branchResult_predictFail <= 1'b0;
      queue_2_exceptionInfo_exception <= 1'b0;
      queue_2_exceptionInfo_eCode <= 6'h00;
      queue_2_exceptionInfo_eSubCode <= 1'b0;
      queue_2_pc <= 32'h00000000;
      queue_2_prd <= 6'h00;
      queue_2_psrc_0 <= 6'h00;
      queue_2_psrc_1 <= 6'h00;
      queue_2_imm <= 32'h00000000;
      queue_2_uop_divuOp <= DIVUOp_div;
      queue_2_srcReady_0 <= 1'b0;
      queue_2_srcReady_1 <= 1'b0;
      queue_3_valid <= 1'b0;
      queue_3_robIdx <= 5'h00;
      queue_3_branchResult_targetPC <= 32'h00000000;
      queue_3_branchResult_branchResult <= 1'b0;
      queue_3_branchResult_predictFail <= 1'b0;
      queue_3_exceptionInfo_exception <= 1'b0;
      queue_3_exceptionInfo_eCode <= 6'h00;
      queue_3_exceptionInfo_eSubCode <= 1'b0;
      queue_3_pc <= 32'h00000000;
      queue_3_prd <= 6'h00;
      queue_3_psrc_0 <= 6'h00;
      queue_3_psrc_1 <= 6'h00;
      queue_3_imm <= 32'h00000000;
      queue_3_uop_divuOp <= DIVUOp_div;
      queue_3_srcReady_0 <= 1'b0;
      queue_3_srcReady_1 <= 1'b0;
    end else begin
      queue_0_valid <= queueNext_0_valid;
      queue_0_robIdx <= queueNext_0_robIdx;
      queue_0_branchResult_targetPC <= queueNext_0_branchResult_targetPC;
      queue_0_branchResult_branchResult <= queueNext_0_branchResult_branchResult;
      queue_0_branchResult_predictFail <= queueNext_0_branchResult_predictFail;
      queue_0_exceptionInfo_exception <= queueNext_0_exceptionInfo_exception;
      queue_0_exceptionInfo_eCode <= queueNext_0_exceptionInfo_eCode;
      queue_0_exceptionInfo_eSubCode <= queueNext_0_exceptionInfo_eSubCode;
      queue_0_pc <= queueNext_0_pc;
      queue_0_prd <= queueNext_0_prd;
      queue_0_psrc_0 <= queueNext_0_psrc_0;
      queue_0_psrc_1 <= queueNext_0_psrc_1;
      queue_0_imm <= queueNext_0_imm;
      queue_0_uop_divuOp <= queueNext_0_uop_divuOp;
      queue_0_srcReady_0 <= queueNext_0_srcReady_0;
      queue_0_srcReady_1 <= queueNext_0_srcReady_1;
      queue_1_valid <= queueNext_1_valid;
      queue_1_robIdx <= queueNext_1_robIdx;
      queue_1_branchResult_targetPC <= queueNext_1_branchResult_targetPC;
      queue_1_branchResult_branchResult <= queueNext_1_branchResult_branchResult;
      queue_1_branchResult_predictFail <= queueNext_1_branchResult_predictFail;
      queue_1_exceptionInfo_exception <= queueNext_1_exceptionInfo_exception;
      queue_1_exceptionInfo_eCode <= queueNext_1_exceptionInfo_eCode;
      queue_1_exceptionInfo_eSubCode <= queueNext_1_exceptionInfo_eSubCode;
      queue_1_pc <= queueNext_1_pc;
      queue_1_prd <= queueNext_1_prd;
      queue_1_psrc_0 <= queueNext_1_psrc_0;
      queue_1_psrc_1 <= queueNext_1_psrc_1;
      queue_1_imm <= queueNext_1_imm;
      queue_1_uop_divuOp <= queueNext_1_uop_divuOp;
      queue_1_srcReady_0 <= queueNext_1_srcReady_0;
      queue_1_srcReady_1 <= queueNext_1_srcReady_1;
      queue_2_valid <= queueNext_2_valid;
      queue_2_robIdx <= queueNext_2_robIdx;
      queue_2_branchResult_targetPC <= queueNext_2_branchResult_targetPC;
      queue_2_branchResult_branchResult <= queueNext_2_branchResult_branchResult;
      queue_2_branchResult_predictFail <= queueNext_2_branchResult_predictFail;
      queue_2_exceptionInfo_exception <= queueNext_2_exceptionInfo_exception;
      queue_2_exceptionInfo_eCode <= queueNext_2_exceptionInfo_eCode;
      queue_2_exceptionInfo_eSubCode <= queueNext_2_exceptionInfo_eSubCode;
      queue_2_pc <= queueNext_2_pc;
      queue_2_prd <= queueNext_2_prd;
      queue_2_psrc_0 <= queueNext_2_psrc_0;
      queue_2_psrc_1 <= queueNext_2_psrc_1;
      queue_2_imm <= queueNext_2_imm;
      queue_2_uop_divuOp <= queueNext_2_uop_divuOp;
      queue_2_srcReady_0 <= queueNext_2_srcReady_0;
      queue_2_srcReady_1 <= queueNext_2_srcReady_1;
      queue_3_valid <= queueNext_3_valid;
      queue_3_robIdx <= queueNext_3_robIdx;
      queue_3_branchResult_targetPC <= queueNext_3_branchResult_targetPC;
      queue_3_branchResult_branchResult <= queueNext_3_branchResult_branchResult;
      queue_3_branchResult_predictFail <= queueNext_3_branchResult_predictFail;
      queue_3_exceptionInfo_exception <= queueNext_3_exceptionInfo_exception;
      queue_3_exceptionInfo_eCode <= queueNext_3_exceptionInfo_eCode;
      queue_3_exceptionInfo_eSubCode <= queueNext_3_exceptionInfo_eSubCode;
      queue_3_pc <= queueNext_3_pc;
      queue_3_prd <= queueNext_3_prd;
      queue_3_psrc_0 <= queueNext_3_psrc_0;
      queue_3_psrc_1 <= queueNext_3_psrc_1;
      queue_3_imm <= queueNext_3_imm;
      queue_3_uop_divuOp <= queueNext_3_uop_divuOp;
      queue_3_srcReady_0 <= queueNext_3_srcReady_0;
      queue_3_srcReady_1 <= queueNext_3_srcReady_1;
    end
  end


endmodule

module IssueQueue_2 (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [4:0]    io_input_payload_robIdx,
  input  wire [31:0]   io_input_payload_branchResult_targetPC,
  input  wire          io_input_payload_branchResult_branchResult,
  input  wire          io_input_payload_branchResult_predictFail,
  input  wire          io_input_payload_exceptionInfo_exception,
  input  wire [5:0]    io_input_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_input_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_payload_pc,
  input  wire [5:0]    io_input_payload_prd,
  input  wire [5:0]    io_input_payload_psrc_0,
  input  wire [5:0]    io_input_payload_psrc_1,
  input  wire [31:0]   io_input_payload_imm,
  input  wire [1:0]    io_input_payload_uop_muluOp,
  input  wire          io_input_payload_srcReady_0,
  input  wire          io_input_payload_srcReady_1,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [4:0]    io_output_payload_robIdx,
  output wire [31:0]   io_output_payload_branchResult_targetPC,
  output wire          io_output_payload_branchResult_branchResult,
  output wire          io_output_payload_branchResult_predictFail,
  output wire          io_output_payload_exceptionInfo_exception,
  output wire [5:0]    io_output_payload_exceptionInfo_eCode,
  output wire [0:0]    io_output_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_output_payload_pc,
  output wire [5:0]    io_output_payload_prd,
  output wire [5:0]    io_output_payload_psrc_0,
  output wire [5:0]    io_output_payload_psrc_1,
  output wire [31:0]   io_output_payload_imm,
  output wire [1:0]    io_output_payload_uop_muluOp,
  input  wire [5:0]    io_writebackSignal_0,
  input  wire [5:0]    io_writebackSignal_1,
  input  wire [5:0]    io_writebackSignal_2,
  input  wire [5:0]    io_writebackSignal_3,
  input  wire [5:0]    io_writebackSignal_4,
  input  wire          io_earlyWakeup_0_valid,
  input  wire [5:0]    io_earlyWakeup_0_payload,
  input  wire          io_earlyWakeup_1_valid,
  input  wire [5:0]    io_earlyWakeup_1_payload,
  input  wire          aclk,
  input  wire          cpuClockingArea_areaFlushReset_newReset
);
  localparam MULUOp_mullo = 2'd0;
  localparam MULUOp_mulhi = 2'd1;
  localparam MULUOp_mulhiu = 2'd2;

  wire       [3:0]    _zz_readyToIssue_ohFirst_masked;
  wire       [4:0]    _zz_emptyEntry_ohFirst_masked;
  wire                _zz_appendEntry_srcReady_0;
  wire       [0:0]    _zz_appendEntry_srcReady_0_1;
  wire       [0:0]    _zz_appendEntry_srcReady_0_2;
  wire                _zz_appendEntry_srcReady_1;
  wire       [0:0]    _zz_appendEntry_srcReady_1_1;
  wire       [0:0]    _zz_appendEntry_srcReady_1_2;
  wire                _zz_updatedEntry_0_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_0_2;
  wire                _zz_updatedEntry_0_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_1_2;
  wire                _zz_updatedEntry_1_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_0_2;
  wire                _zz_updatedEntry_1_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_1_2;
  wire                _zz_updatedEntry_2_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_0_2;
  wire                _zz_updatedEntry_2_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_1_2;
  wire                _zz_updatedEntry_3_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_0_2;
  wire                _zz_updatedEntry_3_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_1_2;
  reg                 _zz_issueEntry_valid_4;
  reg        [4:0]    _zz_issueEntry_robIdx;
  reg        [31:0]   _zz_issueEntry_branchResult_targetPC;
  reg                 _zz_issueEntry_branchResult_branchResult;
  reg                 _zz_issueEntry_branchResult_predictFail;
  reg                 _zz_issueEntry_exceptionInfo_exception;
  reg        [5:0]    _zz_issueEntry_exceptionInfo_eCode;
  reg        [0:0]    _zz_issueEntry_exceptionInfo_eSubCode;
  reg        [31:0]   _zz_issueEntry_pc;
  reg        [5:0]    _zz_issueEntry_prd;
  reg        [5:0]    _zz_issueEntry_psrc_0;
  reg        [5:0]    _zz_issueEntry_psrc_1;
  reg        [31:0]   _zz_issueEntry_imm;
  reg        [1:0]    _zz_issueEntry_uop_muluOp;
  reg                 _zz_issueEntry_srcReady_0;
  reg                 _zz_issueEntry_srcReady_1;
  reg                 queue_0_valid;
  reg        [4:0]    queue_0_robIdx;
  reg        [31:0]   queue_0_branchResult_targetPC;
  reg                 queue_0_branchResult_branchResult;
  reg                 queue_0_branchResult_predictFail;
  reg                 queue_0_exceptionInfo_exception;
  reg        [5:0]    queue_0_exceptionInfo_eCode;
  reg        [0:0]    queue_0_exceptionInfo_eSubCode;
  reg        [31:0]   queue_0_pc;
  reg        [5:0]    queue_0_prd;
  reg        [5:0]    queue_0_psrc_0;
  reg        [5:0]    queue_0_psrc_1;
  reg        [31:0]   queue_0_imm;
  reg        [1:0]    queue_0_uop_muluOp;
  reg                 queue_0_srcReady_0;
  reg                 queue_0_srcReady_1;
  reg                 queue_1_valid;
  reg        [4:0]    queue_1_robIdx;
  reg        [31:0]   queue_1_branchResult_targetPC;
  reg                 queue_1_branchResult_branchResult;
  reg                 queue_1_branchResult_predictFail;
  reg                 queue_1_exceptionInfo_exception;
  reg        [5:0]    queue_1_exceptionInfo_eCode;
  reg        [0:0]    queue_1_exceptionInfo_eSubCode;
  reg        [31:0]   queue_1_pc;
  reg        [5:0]    queue_1_prd;
  reg        [5:0]    queue_1_psrc_0;
  reg        [5:0]    queue_1_psrc_1;
  reg        [31:0]   queue_1_imm;
  reg        [1:0]    queue_1_uop_muluOp;
  reg                 queue_1_srcReady_0;
  reg                 queue_1_srcReady_1;
  reg                 queue_2_valid;
  reg        [4:0]    queue_2_robIdx;
  reg        [31:0]   queue_2_branchResult_targetPC;
  reg                 queue_2_branchResult_branchResult;
  reg                 queue_2_branchResult_predictFail;
  reg                 queue_2_exceptionInfo_exception;
  reg        [5:0]    queue_2_exceptionInfo_eCode;
  reg        [0:0]    queue_2_exceptionInfo_eSubCode;
  reg        [31:0]   queue_2_pc;
  reg        [5:0]    queue_2_prd;
  reg        [5:0]    queue_2_psrc_0;
  reg        [5:0]    queue_2_psrc_1;
  reg        [31:0]   queue_2_imm;
  reg        [1:0]    queue_2_uop_muluOp;
  reg                 queue_2_srcReady_0;
  reg                 queue_2_srcReady_1;
  reg                 queue_3_valid;
  reg        [4:0]    queue_3_robIdx;
  reg        [31:0]   queue_3_branchResult_targetPC;
  reg                 queue_3_branchResult_branchResult;
  reg                 queue_3_branchResult_predictFail;
  reg                 queue_3_exceptionInfo_exception;
  reg        [5:0]    queue_3_exceptionInfo_eCode;
  reg        [0:0]    queue_3_exceptionInfo_eSubCode;
  reg        [31:0]   queue_3_pc;
  reg        [5:0]    queue_3_prd;
  reg        [5:0]    queue_3_psrc_0;
  reg        [5:0]    queue_3_psrc_1;
  reg        [31:0]   queue_3_imm;
  reg        [1:0]    queue_3_uop_muluOp;
  reg                 queue_3_srcReady_0;
  reg                 queue_3_srcReady_1;
  reg        [3:0]    readyToIssue;
  wire       [3:0]    readyToIssue_ohFirst_input;
  wire       [3:0]    readyToIssue_ohFirst_masked;
  wire       [3:0]    issueVector;
  reg        [3:0]    shiftAhead;
  reg        [4:0]    emptyEntry;
  wire       [4:0]    emptyEntry_ohFirst_input;
  wire       [4:0]    emptyEntry_ohFirst_masked;
  wire       [4:0]    writeVector;
  wire                updatedEntry_0_valid;
  wire       [4:0]    updatedEntry_0_robIdx;
  wire       [31:0]   updatedEntry_0_branchResult_targetPC;
  wire                updatedEntry_0_branchResult_branchResult;
  wire                updatedEntry_0_branchResult_predictFail;
  wire                updatedEntry_0_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_0_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_0_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_0_pc;
  wire       [5:0]    updatedEntry_0_prd;
  wire       [5:0]    updatedEntry_0_psrc_0;
  wire       [5:0]    updatedEntry_0_psrc_1;
  wire       [31:0]   updatedEntry_0_imm;
  wire       [1:0]    updatedEntry_0_uop_muluOp;
  reg                 updatedEntry_0_srcReady_0;
  reg                 updatedEntry_0_srcReady_1;
  wire                updatedEntry_1_valid;
  wire       [4:0]    updatedEntry_1_robIdx;
  wire       [31:0]   updatedEntry_1_branchResult_targetPC;
  wire                updatedEntry_1_branchResult_branchResult;
  wire                updatedEntry_1_branchResult_predictFail;
  wire                updatedEntry_1_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_1_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_1_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_1_pc;
  wire       [5:0]    updatedEntry_1_prd;
  wire       [5:0]    updatedEntry_1_psrc_0;
  wire       [5:0]    updatedEntry_1_psrc_1;
  wire       [31:0]   updatedEntry_1_imm;
  wire       [1:0]    updatedEntry_1_uop_muluOp;
  reg                 updatedEntry_1_srcReady_0;
  reg                 updatedEntry_1_srcReady_1;
  wire                updatedEntry_2_valid;
  wire       [4:0]    updatedEntry_2_robIdx;
  wire       [31:0]   updatedEntry_2_branchResult_targetPC;
  wire                updatedEntry_2_branchResult_branchResult;
  wire                updatedEntry_2_branchResult_predictFail;
  wire                updatedEntry_2_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_2_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_2_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_2_pc;
  wire       [5:0]    updatedEntry_2_prd;
  wire       [5:0]    updatedEntry_2_psrc_0;
  wire       [5:0]    updatedEntry_2_psrc_1;
  wire       [31:0]   updatedEntry_2_imm;
  wire       [1:0]    updatedEntry_2_uop_muluOp;
  reg                 updatedEntry_2_srcReady_0;
  reg                 updatedEntry_2_srcReady_1;
  wire                updatedEntry_3_valid;
  wire       [4:0]    updatedEntry_3_robIdx;
  wire       [31:0]   updatedEntry_3_branchResult_targetPC;
  wire                updatedEntry_3_branchResult_branchResult;
  wire                updatedEntry_3_branchResult_predictFail;
  wire                updatedEntry_3_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_3_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_3_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_3_pc;
  wire       [5:0]    updatedEntry_3_prd;
  wire       [5:0]    updatedEntry_3_psrc_0;
  wire       [5:0]    updatedEntry_3_psrc_1;
  wire       [31:0]   updatedEntry_3_imm;
  wire       [1:0]    updatedEntry_3_uop_muluOp;
  reg                 updatedEntry_3_srcReady_0;
  reg                 updatedEntry_3_srcReady_1;
  wire                appendEntry_valid;
  wire       [4:0]    appendEntry_robIdx;
  wire       [31:0]   appendEntry_branchResult_targetPC;
  wire                appendEntry_branchResult_branchResult;
  wire                appendEntry_branchResult_predictFail;
  wire                appendEntry_exceptionInfo_exception;
  wire       [5:0]    appendEntry_exceptionInfo_eCode;
  wire       [0:0]    appendEntry_exceptionInfo_eSubCode;
  wire       [31:0]   appendEntry_pc;
  wire       [5:0]    appendEntry_prd;
  wire       [5:0]    appendEntry_psrc_0;
  wire       [5:0]    appendEntry_psrc_1;
  wire       [31:0]   appendEntry_imm;
  wire       [1:0]    appendEntry_uop_muluOp;
  wire                appendEntry_srcReady_0;
  wire                appendEntry_srcReady_1;
  reg                 queueNext_0_valid;
  reg        [4:0]    queueNext_0_robIdx;
  reg        [31:0]   queueNext_0_branchResult_targetPC;
  reg                 queueNext_0_branchResult_branchResult;
  reg                 queueNext_0_branchResult_predictFail;
  reg                 queueNext_0_exceptionInfo_exception;
  reg        [5:0]    queueNext_0_exceptionInfo_eCode;
  reg        [0:0]    queueNext_0_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_0_pc;
  reg        [5:0]    queueNext_0_prd;
  reg        [5:0]    queueNext_0_psrc_0;
  reg        [5:0]    queueNext_0_psrc_1;
  reg        [31:0]   queueNext_0_imm;
  reg        [1:0]    queueNext_0_uop_muluOp;
  reg                 queueNext_0_srcReady_0;
  reg                 queueNext_0_srcReady_1;
  reg                 queueNext_1_valid;
  reg        [4:0]    queueNext_1_robIdx;
  reg        [31:0]   queueNext_1_branchResult_targetPC;
  reg                 queueNext_1_branchResult_branchResult;
  reg                 queueNext_1_branchResult_predictFail;
  reg                 queueNext_1_exceptionInfo_exception;
  reg        [5:0]    queueNext_1_exceptionInfo_eCode;
  reg        [0:0]    queueNext_1_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_1_pc;
  reg        [5:0]    queueNext_1_prd;
  reg        [5:0]    queueNext_1_psrc_0;
  reg        [5:0]    queueNext_1_psrc_1;
  reg        [31:0]   queueNext_1_imm;
  reg        [1:0]    queueNext_1_uop_muluOp;
  reg                 queueNext_1_srcReady_0;
  reg                 queueNext_1_srcReady_1;
  reg                 queueNext_2_valid;
  reg        [4:0]    queueNext_2_robIdx;
  reg        [31:0]   queueNext_2_branchResult_targetPC;
  reg                 queueNext_2_branchResult_branchResult;
  reg                 queueNext_2_branchResult_predictFail;
  reg                 queueNext_2_exceptionInfo_exception;
  reg        [5:0]    queueNext_2_exceptionInfo_eCode;
  reg        [0:0]    queueNext_2_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_2_pc;
  reg        [5:0]    queueNext_2_prd;
  reg        [5:0]    queueNext_2_psrc_0;
  reg        [5:0]    queueNext_2_psrc_1;
  reg        [31:0]   queueNext_2_imm;
  reg        [1:0]    queueNext_2_uop_muluOp;
  reg                 queueNext_2_srcReady_0;
  reg                 queueNext_2_srcReady_1;
  reg                 queueNext_3_valid;
  reg        [4:0]    queueNext_3_robIdx;
  reg        [31:0]   queueNext_3_branchResult_targetPC;
  reg                 queueNext_3_branchResult_branchResult;
  reg                 queueNext_3_branchResult_predictFail;
  reg                 queueNext_3_exceptionInfo_exception;
  reg        [5:0]    queueNext_3_exceptionInfo_eCode;
  reg        [0:0]    queueNext_3_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_3_pc;
  reg        [5:0]    queueNext_3_prd;
  reg        [5:0]    queueNext_3_psrc_0;
  reg        [5:0]    queueNext_3_psrc_1;
  reg        [31:0]   queueNext_3_imm;
  reg        [1:0]    queueNext_3_uop_muluOp;
  reg                 queueNext_3_srcReady_0;
  reg                 queueNext_3_srcReady_1;
  wire                when_IssueQueue_l81;
  wire                when_IssueQueue_l83;
  wire                when_IssueQueue_l96;
  wire                when_IssueQueue_l81_1;
  wire                when_IssueQueue_l83_1;
  wire                when_IssueQueue_l96_1;
  wire                when_IssueQueue_l81_2;
  wire                when_IssueQueue_l83_2;
  wire                when_IssueQueue_l96_2;
  wire                when_IssueQueue_l81_3;
  wire                when_IssueQueue_l89;
  wire                when_IssueQueue_l96_3;
  wire                io_output_fire;
  wire                _zz_issueEntry_valid;
  wire                _zz_issueEntry_valid_1;
  wire                _zz_issueEntry_valid_2;
  wire       [1:0]    _zz_issueEntry_valid_3;
  wire                issueEntry_valid;
  wire       [4:0]    issueEntry_robIdx;
  wire       [31:0]   issueEntry_branchResult_targetPC;
  wire                issueEntry_branchResult_branchResult;
  wire                issueEntry_branchResult_predictFail;
  wire                issueEntry_exceptionInfo_exception;
  wire       [5:0]    issueEntry_exceptionInfo_eCode;
  wire       [0:0]    issueEntry_exceptionInfo_eSubCode;
  wire       [31:0]   issueEntry_pc;
  wire       [5:0]    issueEntry_prd;
  wire       [5:0]    issueEntry_psrc_0;
  wire       [5:0]    issueEntry_psrc_1;
  wire       [31:0]   issueEntry_imm;
  wire       [1:0]    issueEntry_uop_muluOp;
  wire                issueEntry_srcReady_0;
  wire                issueEntry_srcReady_1;
  `ifndef SYNTHESIS
  reg [47:0] io_input_payload_uop_muluOp_string;
  reg [47:0] io_output_payload_uop_muluOp_string;
  reg [47:0] queue_0_uop_muluOp_string;
  reg [47:0] queue_1_uop_muluOp_string;
  reg [47:0] queue_2_uop_muluOp_string;
  reg [47:0] queue_3_uop_muluOp_string;
  reg [47:0] updatedEntry_0_uop_muluOp_string;
  reg [47:0] updatedEntry_1_uop_muluOp_string;
  reg [47:0] updatedEntry_2_uop_muluOp_string;
  reg [47:0] updatedEntry_3_uop_muluOp_string;
  reg [47:0] appendEntry_uop_muluOp_string;
  reg [47:0] queueNext_0_uop_muluOp_string;
  reg [47:0] queueNext_1_uop_muluOp_string;
  reg [47:0] queueNext_2_uop_muluOp_string;
  reg [47:0] queueNext_3_uop_muluOp_string;
  reg [47:0] issueEntry_uop_muluOp_string;
  `endif


  assign _zz_readyToIssue_ohFirst_masked = (readyToIssue_ohFirst_input - 4'b0001);
  assign _zz_emptyEntry_ohFirst_masked = (emptyEntry_ohFirst_input - 5'h01);
  assign _zz_appendEntry_srcReady_0 = (io_input_payload_psrc_0 == io_writebackSignal_2);
  assign _zz_appendEntry_srcReady_0_1 = (io_input_payload_psrc_0 == io_writebackSignal_1);
  assign _zz_appendEntry_srcReady_0_2 = (io_input_payload_psrc_0 == io_writebackSignal_0);
  assign _zz_appendEntry_srcReady_1 = (io_input_payload_psrc_1 == io_writebackSignal_2);
  assign _zz_appendEntry_srcReady_1_1 = (io_input_payload_psrc_1 == io_writebackSignal_1);
  assign _zz_appendEntry_srcReady_1_2 = (io_input_payload_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_0_srcReady_0 = (queue_0_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_0_srcReady_0_1 = (queue_0_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_0_srcReady_0_2 = (queue_0_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_0_srcReady_1 = (queue_0_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_0_srcReady_1_1 = (queue_0_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_0_srcReady_1_2 = (queue_0_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_1_srcReady_0 = (queue_1_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_1_srcReady_0_1 = (queue_1_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_1_srcReady_0_2 = (queue_1_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_1_srcReady_1 = (queue_1_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_1_srcReady_1_1 = (queue_1_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_1_srcReady_1_2 = (queue_1_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_2_srcReady_0 = (queue_2_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_2_srcReady_0_1 = (queue_2_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_2_srcReady_0_2 = (queue_2_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_2_srcReady_1 = (queue_2_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_2_srcReady_1_1 = (queue_2_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_2_srcReady_1_2 = (queue_2_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_3_srcReady_0 = (queue_3_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_3_srcReady_0_1 = (queue_3_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_3_srcReady_0_2 = (queue_3_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_3_srcReady_1 = (queue_3_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_3_srcReady_1_1 = (queue_3_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_3_srcReady_1_2 = (queue_3_psrc_1 == io_writebackSignal_0);
  always @(*) begin
    case(_zz_issueEntry_valid_3)
      2'b00 : begin
        _zz_issueEntry_valid_4 = queue_0_valid;
        _zz_issueEntry_robIdx = queue_0_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_0_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_0_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_0_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_0_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_0_pc;
        _zz_issueEntry_prd = queue_0_prd;
        _zz_issueEntry_psrc_0 = queue_0_psrc_0;
        _zz_issueEntry_psrc_1 = queue_0_psrc_1;
        _zz_issueEntry_imm = queue_0_imm;
        _zz_issueEntry_uop_muluOp = queue_0_uop_muluOp;
        _zz_issueEntry_srcReady_0 = queue_0_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_0_srcReady_1;
      end
      2'b01 : begin
        _zz_issueEntry_valid_4 = queue_1_valid;
        _zz_issueEntry_robIdx = queue_1_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_1_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_1_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_1_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_1_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_1_pc;
        _zz_issueEntry_prd = queue_1_prd;
        _zz_issueEntry_psrc_0 = queue_1_psrc_0;
        _zz_issueEntry_psrc_1 = queue_1_psrc_1;
        _zz_issueEntry_imm = queue_1_imm;
        _zz_issueEntry_uop_muluOp = queue_1_uop_muluOp;
        _zz_issueEntry_srcReady_0 = queue_1_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_1_srcReady_1;
      end
      2'b10 : begin
        _zz_issueEntry_valid_4 = queue_2_valid;
        _zz_issueEntry_robIdx = queue_2_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_2_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_2_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_2_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_2_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_2_pc;
        _zz_issueEntry_prd = queue_2_prd;
        _zz_issueEntry_psrc_0 = queue_2_psrc_0;
        _zz_issueEntry_psrc_1 = queue_2_psrc_1;
        _zz_issueEntry_imm = queue_2_imm;
        _zz_issueEntry_uop_muluOp = queue_2_uop_muluOp;
        _zz_issueEntry_srcReady_0 = queue_2_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_2_srcReady_1;
      end
      default : begin
        _zz_issueEntry_valid_4 = queue_3_valid;
        _zz_issueEntry_robIdx = queue_3_robIdx;
        _zz_issueEntry_branchResult_targetPC = queue_3_branchResult_targetPC;
        _zz_issueEntry_branchResult_branchResult = queue_3_branchResult_branchResult;
        _zz_issueEntry_branchResult_predictFail = queue_3_branchResult_predictFail;
        _zz_issueEntry_exceptionInfo_exception = queue_3_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_3_pc;
        _zz_issueEntry_prd = queue_3_prd;
        _zz_issueEntry_psrc_0 = queue_3_psrc_0;
        _zz_issueEntry_psrc_1 = queue_3_psrc_1;
        _zz_issueEntry_imm = queue_3_imm;
        _zz_issueEntry_uop_muluOp = queue_3_uop_muluOp;
        _zz_issueEntry_srcReady_0 = queue_3_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_3_srcReady_1;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_uop_muluOp)
      MULUOp_mullo : io_input_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : io_input_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : io_input_payload_uop_muluOp_string = "mulhiu";
      default : io_input_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_uop_muluOp)
      MULUOp_mullo : io_output_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : io_output_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : io_output_payload_uop_muluOp_string = "mulhiu";
      default : io_output_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queue_0_uop_muluOp)
      MULUOp_mullo : queue_0_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : queue_0_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : queue_0_uop_muluOp_string = "mulhiu";
      default : queue_0_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queue_1_uop_muluOp)
      MULUOp_mullo : queue_1_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : queue_1_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : queue_1_uop_muluOp_string = "mulhiu";
      default : queue_1_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queue_2_uop_muluOp)
      MULUOp_mullo : queue_2_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : queue_2_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : queue_2_uop_muluOp_string = "mulhiu";
      default : queue_2_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queue_3_uop_muluOp)
      MULUOp_mullo : queue_3_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : queue_3_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : queue_3_uop_muluOp_string = "mulhiu";
      default : queue_3_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_uop_muluOp)
      MULUOp_mullo : updatedEntry_0_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : updatedEntry_0_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : updatedEntry_0_uop_muluOp_string = "mulhiu";
      default : updatedEntry_0_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_uop_muluOp)
      MULUOp_mullo : updatedEntry_1_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : updatedEntry_1_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : updatedEntry_1_uop_muluOp_string = "mulhiu";
      default : updatedEntry_1_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_uop_muluOp)
      MULUOp_mullo : updatedEntry_2_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : updatedEntry_2_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : updatedEntry_2_uop_muluOp_string = "mulhiu";
      default : updatedEntry_2_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_uop_muluOp)
      MULUOp_mullo : updatedEntry_3_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : updatedEntry_3_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : updatedEntry_3_uop_muluOp_string = "mulhiu";
      default : updatedEntry_3_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(appendEntry_uop_muluOp)
      MULUOp_mullo : appendEntry_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : appendEntry_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : appendEntry_uop_muluOp_string = "mulhiu";
      default : appendEntry_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queueNext_0_uop_muluOp)
      MULUOp_mullo : queueNext_0_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : queueNext_0_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : queueNext_0_uop_muluOp_string = "mulhiu";
      default : queueNext_0_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queueNext_1_uop_muluOp)
      MULUOp_mullo : queueNext_1_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : queueNext_1_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : queueNext_1_uop_muluOp_string = "mulhiu";
      default : queueNext_1_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queueNext_2_uop_muluOp)
      MULUOp_mullo : queueNext_2_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : queueNext_2_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : queueNext_2_uop_muluOp_string = "mulhiu";
      default : queueNext_2_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(queueNext_3_uop_muluOp)
      MULUOp_mullo : queueNext_3_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : queueNext_3_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : queueNext_3_uop_muluOp_string = "mulhiu";
      default : queueNext_3_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(issueEntry_uop_muluOp)
      MULUOp_mullo : issueEntry_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : issueEntry_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : issueEntry_uop_muluOp_string = "mulhiu";
      default : issueEntry_uop_muluOp_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    readyToIssue[0] = ((queue_0_valid && queue_0_srcReady_0) && queue_0_srcReady_1);
    readyToIssue[1] = ((queue_1_valid && queue_1_srcReady_0) && queue_1_srcReady_1);
    readyToIssue[2] = ((queue_2_valid && queue_2_srcReady_0) && queue_2_srcReady_1);
    readyToIssue[3] = ((queue_3_valid && queue_3_srcReady_0) && queue_3_srcReady_1);
  end

  assign readyToIssue_ohFirst_input = readyToIssue;
  assign readyToIssue_ohFirst_masked = (readyToIssue_ohFirst_input & (~ _zz_readyToIssue_ohFirst_masked));
  assign issueVector = readyToIssue_ohFirst_masked;
  always @(*) begin
    emptyEntry[0] = (! queue_0_valid);
    emptyEntry[1] = (! queue_1_valid);
    emptyEntry[2] = (! queue_2_valid);
    emptyEntry[3] = (! queue_3_valid);
    emptyEntry[4] = 1'b1;
    emptyEntry[0] = (! queue_0_valid);
    emptyEntry[1] = (! queue_1_valid);
    emptyEntry[2] = (! queue_2_valid);
    emptyEntry[3] = (! queue_3_valid);
  end

  assign emptyEntry_ohFirst_input = emptyEntry;
  assign emptyEntry_ohFirst_masked = (emptyEntry_ohFirst_input & (~ _zz_emptyEntry_ohFirst_masked));
  assign writeVector = emptyEntry_ohFirst_masked;
  assign appendEntry_valid = io_input_valid;
  assign appendEntry_robIdx = io_input_payload_robIdx;
  assign appendEntry_branchResult_targetPC = io_input_payload_branchResult_targetPC;
  assign appendEntry_branchResult_branchResult = io_input_payload_branchResult_branchResult;
  assign appendEntry_branchResult_predictFail = io_input_payload_branchResult_predictFail;
  assign appendEntry_exceptionInfo_exception = io_input_payload_exceptionInfo_exception;
  assign appendEntry_exceptionInfo_eCode = io_input_payload_exceptionInfo_eCode;
  assign appendEntry_exceptionInfo_eSubCode = io_input_payload_exceptionInfo_eSubCode;
  assign appendEntry_pc = io_input_payload_pc;
  assign appendEntry_prd = io_input_payload_prd;
  assign appendEntry_psrc_0 = io_input_payload_psrc_0;
  assign appendEntry_psrc_1 = io_input_payload_psrc_1;
  assign appendEntry_imm = io_input_payload_imm;
  assign appendEntry_uop_muluOp = io_input_payload_uop_muluOp;
  assign appendEntry_srcReady_0 = ((io_input_payload_srcReady_0 || (|{(io_input_payload_psrc_0 == io_writebackSignal_4),{(io_input_payload_psrc_0 == io_writebackSignal_3),{_zz_appendEntry_srcReady_0,{_zz_appendEntry_srcReady_0_1,_zz_appendEntry_srcReady_0_2}}}})) || (|{((io_input_payload_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((io_input_payload_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}));
  assign appendEntry_srcReady_1 = ((io_input_payload_srcReady_1 || (|{(io_input_payload_psrc_1 == io_writebackSignal_4),{(io_input_payload_psrc_1 == io_writebackSignal_3),{_zz_appendEntry_srcReady_1,{_zz_appendEntry_srcReady_1_1,_zz_appendEntry_srcReady_1_2}}}})) || (|{((io_input_payload_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((io_input_payload_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}));
  assign updatedEntry_0_valid = queue_0_valid;
  assign updatedEntry_0_robIdx = queue_0_robIdx;
  assign updatedEntry_0_branchResult_targetPC = queue_0_branchResult_targetPC;
  assign updatedEntry_0_branchResult_branchResult = queue_0_branchResult_branchResult;
  assign updatedEntry_0_branchResult_predictFail = queue_0_branchResult_predictFail;
  assign updatedEntry_0_exceptionInfo_exception = queue_0_exceptionInfo_exception;
  assign updatedEntry_0_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
  assign updatedEntry_0_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
  assign updatedEntry_0_pc = queue_0_pc;
  assign updatedEntry_0_prd = queue_0_prd;
  assign updatedEntry_0_psrc_0 = queue_0_psrc_0;
  assign updatedEntry_0_psrc_1 = queue_0_psrc_1;
  assign updatedEntry_0_imm = queue_0_imm;
  assign updatedEntry_0_uop_muluOp = queue_0_uop_muluOp;
  always @(*) begin
    updatedEntry_0_srcReady_0 = queue_0_srcReady_0;
    updatedEntry_0_srcReady_0 = ((queue_0_srcReady_0 || (|{(queue_0_psrc_0 == io_writebackSignal_4),{(queue_0_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_0_srcReady_0,{_zz_updatedEntry_0_srcReady_0_1,_zz_updatedEntry_0_srcReady_0_2}}}})) || (|{((queue_0_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_0_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}));
  end

  always @(*) begin
    updatedEntry_0_srcReady_1 = queue_0_srcReady_1;
    updatedEntry_0_srcReady_1 = ((queue_0_srcReady_1 || (|{(queue_0_psrc_1 == io_writebackSignal_4),{(queue_0_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_0_srcReady_1,{_zz_updatedEntry_0_srcReady_1_1,_zz_updatedEntry_0_srcReady_1_2}}}})) || (|{((queue_0_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_0_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}));
  end

  assign updatedEntry_1_valid = queue_1_valid;
  assign updatedEntry_1_robIdx = queue_1_robIdx;
  assign updatedEntry_1_branchResult_targetPC = queue_1_branchResult_targetPC;
  assign updatedEntry_1_branchResult_branchResult = queue_1_branchResult_branchResult;
  assign updatedEntry_1_branchResult_predictFail = queue_1_branchResult_predictFail;
  assign updatedEntry_1_exceptionInfo_exception = queue_1_exceptionInfo_exception;
  assign updatedEntry_1_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
  assign updatedEntry_1_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
  assign updatedEntry_1_pc = queue_1_pc;
  assign updatedEntry_1_prd = queue_1_prd;
  assign updatedEntry_1_psrc_0 = queue_1_psrc_0;
  assign updatedEntry_1_psrc_1 = queue_1_psrc_1;
  assign updatedEntry_1_imm = queue_1_imm;
  assign updatedEntry_1_uop_muluOp = queue_1_uop_muluOp;
  always @(*) begin
    updatedEntry_1_srcReady_0 = queue_1_srcReady_0;
    updatedEntry_1_srcReady_0 = ((queue_1_srcReady_0 || (|{(queue_1_psrc_0 == io_writebackSignal_4),{(queue_1_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_1_srcReady_0,{_zz_updatedEntry_1_srcReady_0_1,_zz_updatedEntry_1_srcReady_0_2}}}})) || (|{((queue_1_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_1_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}));
  end

  always @(*) begin
    updatedEntry_1_srcReady_1 = queue_1_srcReady_1;
    updatedEntry_1_srcReady_1 = ((queue_1_srcReady_1 || (|{(queue_1_psrc_1 == io_writebackSignal_4),{(queue_1_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_1_srcReady_1,{_zz_updatedEntry_1_srcReady_1_1,_zz_updatedEntry_1_srcReady_1_2}}}})) || (|{((queue_1_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_1_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}));
  end

  assign updatedEntry_2_valid = queue_2_valid;
  assign updatedEntry_2_robIdx = queue_2_robIdx;
  assign updatedEntry_2_branchResult_targetPC = queue_2_branchResult_targetPC;
  assign updatedEntry_2_branchResult_branchResult = queue_2_branchResult_branchResult;
  assign updatedEntry_2_branchResult_predictFail = queue_2_branchResult_predictFail;
  assign updatedEntry_2_exceptionInfo_exception = queue_2_exceptionInfo_exception;
  assign updatedEntry_2_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
  assign updatedEntry_2_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
  assign updatedEntry_2_pc = queue_2_pc;
  assign updatedEntry_2_prd = queue_2_prd;
  assign updatedEntry_2_psrc_0 = queue_2_psrc_0;
  assign updatedEntry_2_psrc_1 = queue_2_psrc_1;
  assign updatedEntry_2_imm = queue_2_imm;
  assign updatedEntry_2_uop_muluOp = queue_2_uop_muluOp;
  always @(*) begin
    updatedEntry_2_srcReady_0 = queue_2_srcReady_0;
    updatedEntry_2_srcReady_0 = ((queue_2_srcReady_0 || (|{(queue_2_psrc_0 == io_writebackSignal_4),{(queue_2_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_2_srcReady_0,{_zz_updatedEntry_2_srcReady_0_1,_zz_updatedEntry_2_srcReady_0_2}}}})) || (|{((queue_2_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_2_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}));
  end

  always @(*) begin
    updatedEntry_2_srcReady_1 = queue_2_srcReady_1;
    updatedEntry_2_srcReady_1 = ((queue_2_srcReady_1 || (|{(queue_2_psrc_1 == io_writebackSignal_4),{(queue_2_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_2_srcReady_1,{_zz_updatedEntry_2_srcReady_1_1,_zz_updatedEntry_2_srcReady_1_2}}}})) || (|{((queue_2_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_2_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}));
  end

  assign updatedEntry_3_valid = queue_3_valid;
  assign updatedEntry_3_robIdx = queue_3_robIdx;
  assign updatedEntry_3_branchResult_targetPC = queue_3_branchResult_targetPC;
  assign updatedEntry_3_branchResult_branchResult = queue_3_branchResult_branchResult;
  assign updatedEntry_3_branchResult_predictFail = queue_3_branchResult_predictFail;
  assign updatedEntry_3_exceptionInfo_exception = queue_3_exceptionInfo_exception;
  assign updatedEntry_3_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
  assign updatedEntry_3_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
  assign updatedEntry_3_pc = queue_3_pc;
  assign updatedEntry_3_prd = queue_3_prd;
  assign updatedEntry_3_psrc_0 = queue_3_psrc_0;
  assign updatedEntry_3_psrc_1 = queue_3_psrc_1;
  assign updatedEntry_3_imm = queue_3_imm;
  assign updatedEntry_3_uop_muluOp = queue_3_uop_muluOp;
  always @(*) begin
    updatedEntry_3_srcReady_0 = queue_3_srcReady_0;
    updatedEntry_3_srcReady_0 = ((queue_3_srcReady_0 || (|{(queue_3_psrc_0 == io_writebackSignal_4),{(queue_3_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_3_srcReady_0,{_zz_updatedEntry_3_srcReady_0_1,_zz_updatedEntry_3_srcReady_0_2}}}})) || (|{((queue_3_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_3_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}));
  end

  always @(*) begin
    updatedEntry_3_srcReady_1 = queue_3_srcReady_1;
    updatedEntry_3_srcReady_1 = ((queue_3_srcReady_1 || (|{(queue_3_psrc_1 == io_writebackSignal_4),{(queue_3_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_3_srcReady_1,{_zz_updatedEntry_3_srcReady_1_1,_zz_updatedEntry_3_srcReady_1_2}}}})) || (|{((queue_3_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_3_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}));
  end

  always @(*) begin
    shiftAhead[0] = ((|readyToIssue[0 : 0]) && io_output_ready);
    shiftAhead[1] = ((|readyToIssue[1 : 0]) && io_output_ready);
    shiftAhead[2] = ((|readyToIssue[2 : 0]) && io_output_ready);
    shiftAhead[3] = ((|readyToIssue[3 : 0]) && io_output_ready);
  end

  assign when_IssueQueue_l81 = shiftAhead[0];
  assign when_IssueQueue_l83 = writeVector[1];
  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_valid = appendEntry_valid;
      end else begin
        queueNext_0_valid = queue_1_valid;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_valid = appendEntry_valid;
      end else begin
        queueNext_0_valid = queue_0_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_0_robIdx = queue_1_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_0_robIdx = queue_0_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_0_branchResult_targetPC = queue_1_branchResult_targetPC;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_0_branchResult_targetPC = queue_0_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_0_branchResult_branchResult = queue_1_branchResult_branchResult;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_0_branchResult_branchResult = queue_0_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_0_branchResult_predictFail = queue_1_branchResult_predictFail;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_0_branchResult_predictFail = queue_0_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_0_exceptionInfo_exception = queue_1_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_0_exceptionInfo_exception = queue_0_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_0_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_0_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_0_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_0_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_pc = appendEntry_pc;
      end else begin
        queueNext_0_pc = queue_1_pc;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_pc = appendEntry_pc;
      end else begin
        queueNext_0_pc = queue_0_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_prd = appendEntry_prd;
      end else begin
        queueNext_0_prd = queue_1_prd;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_prd = appendEntry_prd;
      end else begin
        queueNext_0_prd = queue_0_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_0_psrc_0 = queue_1_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_0_psrc_0 = queue_0_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_0_psrc_1 = queue_1_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_0_psrc_1 = queue_0_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_imm = appendEntry_imm;
      end else begin
        queueNext_0_imm = queue_1_imm;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_imm = appendEntry_imm;
      end else begin
        queueNext_0_imm = queue_0_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_uop_muluOp = appendEntry_uop_muluOp;
      end else begin
        queueNext_0_uop_muluOp = queue_1_uop_muluOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_uop_muluOp = appendEntry_uop_muluOp;
      end else begin
        queueNext_0_uop_muluOp = queue_0_uop_muluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_0_srcReady_0 = queue_1_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_0_srcReady_0 = queue_0_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_0_srcReady_1 = queue_1_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_0_srcReady_1 = queue_0_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96 = writeVector[0];
  assign when_IssueQueue_l81_1 = shiftAhead[1];
  assign when_IssueQueue_l83_1 = writeVector[2];
  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_valid = appendEntry_valid;
      end else begin
        queueNext_1_valid = queue_2_valid;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_valid = appendEntry_valid;
      end else begin
        queueNext_1_valid = queue_1_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_1_robIdx = queue_2_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_1_robIdx = queue_1_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_1_branchResult_targetPC = queue_2_branchResult_targetPC;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_1_branchResult_targetPC = queue_1_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_1_branchResult_branchResult = queue_2_branchResult_branchResult;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_1_branchResult_branchResult = queue_1_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_1_branchResult_predictFail = queue_2_branchResult_predictFail;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_1_branchResult_predictFail = queue_1_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_1_exceptionInfo_exception = queue_2_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_1_exceptionInfo_exception = queue_1_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_1_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_1_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_1_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_1_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_pc = appendEntry_pc;
      end else begin
        queueNext_1_pc = queue_2_pc;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_pc = appendEntry_pc;
      end else begin
        queueNext_1_pc = queue_1_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_prd = appendEntry_prd;
      end else begin
        queueNext_1_prd = queue_2_prd;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_prd = appendEntry_prd;
      end else begin
        queueNext_1_prd = queue_1_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_1_psrc_0 = queue_2_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_1_psrc_0 = queue_1_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_1_psrc_1 = queue_2_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_1_psrc_1 = queue_1_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_imm = appendEntry_imm;
      end else begin
        queueNext_1_imm = queue_2_imm;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_imm = appendEntry_imm;
      end else begin
        queueNext_1_imm = queue_1_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_uop_muluOp = appendEntry_uop_muluOp;
      end else begin
        queueNext_1_uop_muluOp = queue_2_uop_muluOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_uop_muluOp = appendEntry_uop_muluOp;
      end else begin
        queueNext_1_uop_muluOp = queue_1_uop_muluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_1_srcReady_0 = queue_2_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_1_srcReady_0 = queue_1_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_1_srcReady_1 = queue_2_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_1_srcReady_1 = queue_1_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_1 = writeVector[1];
  assign when_IssueQueue_l81_2 = shiftAhead[2];
  assign when_IssueQueue_l83_2 = writeVector[3];
  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_valid = appendEntry_valid;
      end else begin
        queueNext_2_valid = queue_3_valid;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_valid = appendEntry_valid;
      end else begin
        queueNext_2_valid = queue_2_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_2_robIdx = queue_3_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_2_robIdx = queue_2_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_2_branchResult_targetPC = queue_3_branchResult_targetPC;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_2_branchResult_targetPC = queue_2_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_2_branchResult_branchResult = queue_3_branchResult_branchResult;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_2_branchResult_branchResult = queue_2_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_2_branchResult_predictFail = queue_3_branchResult_predictFail;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_2_branchResult_predictFail = queue_2_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_2_exceptionInfo_exception = queue_3_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_2_exceptionInfo_exception = queue_2_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_2_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_2_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_2_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_2_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_pc = appendEntry_pc;
      end else begin
        queueNext_2_pc = queue_3_pc;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_pc = appendEntry_pc;
      end else begin
        queueNext_2_pc = queue_2_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_prd = appendEntry_prd;
      end else begin
        queueNext_2_prd = queue_3_prd;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_prd = appendEntry_prd;
      end else begin
        queueNext_2_prd = queue_2_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_2_psrc_0 = queue_3_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_2_psrc_0 = queue_2_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_2_psrc_1 = queue_3_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_2_psrc_1 = queue_2_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_imm = appendEntry_imm;
      end else begin
        queueNext_2_imm = queue_3_imm;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_imm = appendEntry_imm;
      end else begin
        queueNext_2_imm = queue_2_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_uop_muluOp = appendEntry_uop_muluOp;
      end else begin
        queueNext_2_uop_muluOp = queue_3_uop_muluOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_uop_muluOp = appendEntry_uop_muluOp;
      end else begin
        queueNext_2_uop_muluOp = queue_2_uop_muluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_2_srcReady_0 = queue_3_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_2_srcReady_0 = queue_2_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_2_srcReady_1 = queue_3_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_2_srcReady_1 = queue_2_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_2 = writeVector[2];
  assign when_IssueQueue_l81_3 = shiftAhead[3];
  assign when_IssueQueue_l89 = writeVector[4];
  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_valid = appendEntry_valid;
      end else begin
        queueNext_3_valid = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_valid = appendEntry_valid;
      end else begin
        queueNext_3_valid = queue_3_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_3_robIdx = 5'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_3_robIdx = queue_3_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_3_branchResult_targetPC = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchResult_targetPC = appendEntry_branchResult_targetPC;
      end else begin
        queueNext_3_branchResult_targetPC = queue_3_branchResult_targetPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_3_branchResult_branchResult = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchResult_branchResult = appendEntry_branchResult_branchResult;
      end else begin
        queueNext_3_branchResult_branchResult = queue_3_branchResult_branchResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_3_branchResult_predictFail = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchResult_predictFail = appendEntry_branchResult_predictFail;
      end else begin
        queueNext_3_branchResult_predictFail = queue_3_branchResult_predictFail;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_3_exceptionInfo_exception = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_3_exceptionInfo_exception = queue_3_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_3_exceptionInfo_eCode = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_3_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_3_exceptionInfo_eSubCode = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_3_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_pc = appendEntry_pc;
      end else begin
        queueNext_3_pc = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_pc = appendEntry_pc;
      end else begin
        queueNext_3_pc = queue_3_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_prd = appendEntry_prd;
      end else begin
        queueNext_3_prd = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_prd = appendEntry_prd;
      end else begin
        queueNext_3_prd = queue_3_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_3_psrc_0 = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_3_psrc_0 = queue_3_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_3_psrc_1 = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_3_psrc_1 = queue_3_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_imm = appendEntry_imm;
      end else begin
        queueNext_3_imm = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_imm = appendEntry_imm;
      end else begin
        queueNext_3_imm = queue_3_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_uop_muluOp = appendEntry_uop_muluOp;
      end else begin
        queueNext_3_uop_muluOp = MULUOp_mullo;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_uop_muluOp = appendEntry_uop_muluOp;
      end else begin
        queueNext_3_uop_muluOp = queue_3_uop_muluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_3_srcReady_0 = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_3_srcReady_0 = queue_3_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_3_srcReady_1 = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_3_srcReady_1 = queue_3_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_3 = writeVector[3];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_input_ready = ((|emptyEntry[3 : 0]) || io_output_fire);
  assign _zz_issueEntry_valid = issueVector[3];
  assign _zz_issueEntry_valid_1 = (issueVector[1] || _zz_issueEntry_valid);
  assign _zz_issueEntry_valid_2 = (issueVector[2] || _zz_issueEntry_valid);
  assign _zz_issueEntry_valid_3 = {_zz_issueEntry_valid_2,_zz_issueEntry_valid_1};
  assign issueEntry_valid = _zz_issueEntry_valid_4;
  assign issueEntry_robIdx = _zz_issueEntry_robIdx;
  assign issueEntry_branchResult_targetPC = _zz_issueEntry_branchResult_targetPC;
  assign issueEntry_branchResult_branchResult = _zz_issueEntry_branchResult_branchResult;
  assign issueEntry_branchResult_predictFail = _zz_issueEntry_branchResult_predictFail;
  assign issueEntry_exceptionInfo_exception = _zz_issueEntry_exceptionInfo_exception;
  assign issueEntry_exceptionInfo_eCode = _zz_issueEntry_exceptionInfo_eCode;
  assign issueEntry_exceptionInfo_eSubCode = _zz_issueEntry_exceptionInfo_eSubCode;
  assign issueEntry_pc = _zz_issueEntry_pc;
  assign issueEntry_prd = _zz_issueEntry_prd;
  assign issueEntry_psrc_0 = _zz_issueEntry_psrc_0;
  assign issueEntry_psrc_1 = _zz_issueEntry_psrc_1;
  assign issueEntry_imm = _zz_issueEntry_imm;
  assign issueEntry_uop_muluOp = _zz_issueEntry_uop_muluOp;
  assign issueEntry_srcReady_0 = _zz_issueEntry_srcReady_0;
  assign issueEntry_srcReady_1 = _zz_issueEntry_srcReady_1;
  assign io_output_valid = (|readyToIssue);
  assign io_output_payload_robIdx = issueEntry_robIdx;
  assign io_output_payload_branchResult_targetPC = issueEntry_branchResult_targetPC;
  assign io_output_payload_branchResult_branchResult = issueEntry_branchResult_branchResult;
  assign io_output_payload_branchResult_predictFail = issueEntry_branchResult_predictFail;
  assign io_output_payload_exceptionInfo_exception = issueEntry_exceptionInfo_exception;
  assign io_output_payload_exceptionInfo_eCode = issueEntry_exceptionInfo_eCode;
  assign io_output_payload_exceptionInfo_eSubCode = issueEntry_exceptionInfo_eSubCode;
  assign io_output_payload_pc = issueEntry_pc;
  assign io_output_payload_prd = issueEntry_prd;
  assign io_output_payload_psrc_0 = issueEntry_psrc_0;
  assign io_output_payload_psrc_1 = issueEntry_psrc_1;
  assign io_output_payload_imm = issueEntry_imm;
  assign io_output_payload_uop_muluOp = issueEntry_uop_muluOp;
  always @(posedge aclk) begin
    if(!cpuClockingArea_areaFlushReset_newReset) begin
      queue_0_valid <= 1'b0;
      queue_0_robIdx <= 5'h00;
      queue_0_branchResult_targetPC <= 32'h00000000;
      queue_0_branchResult_branchResult <= 1'b0;
      queue_0_branchResult_predictFail <= 1'b0;
      queue_0_exceptionInfo_exception <= 1'b0;
      queue_0_exceptionInfo_eCode <= 6'h00;
      queue_0_exceptionInfo_eSubCode <= 1'b0;
      queue_0_pc <= 32'h00000000;
      queue_0_prd <= 6'h00;
      queue_0_psrc_0 <= 6'h00;
      queue_0_psrc_1 <= 6'h00;
      queue_0_imm <= 32'h00000000;
      queue_0_uop_muluOp <= MULUOp_mullo;
      queue_0_srcReady_0 <= 1'b0;
      queue_0_srcReady_1 <= 1'b0;
      queue_1_valid <= 1'b0;
      queue_1_robIdx <= 5'h00;
      queue_1_branchResult_targetPC <= 32'h00000000;
      queue_1_branchResult_branchResult <= 1'b0;
      queue_1_branchResult_predictFail <= 1'b0;
      queue_1_exceptionInfo_exception <= 1'b0;
      queue_1_exceptionInfo_eCode <= 6'h00;
      queue_1_exceptionInfo_eSubCode <= 1'b0;
      queue_1_pc <= 32'h00000000;
      queue_1_prd <= 6'h00;
      queue_1_psrc_0 <= 6'h00;
      queue_1_psrc_1 <= 6'h00;
      queue_1_imm <= 32'h00000000;
      queue_1_uop_muluOp <= MULUOp_mullo;
      queue_1_srcReady_0 <= 1'b0;
      queue_1_srcReady_1 <= 1'b0;
      queue_2_valid <= 1'b0;
      queue_2_robIdx <= 5'h00;
      queue_2_branchResult_targetPC <= 32'h00000000;
      queue_2_branchResult_branchResult <= 1'b0;
      queue_2_branchResult_predictFail <= 1'b0;
      queue_2_exceptionInfo_exception <= 1'b0;
      queue_2_exceptionInfo_eCode <= 6'h00;
      queue_2_exceptionInfo_eSubCode <= 1'b0;
      queue_2_pc <= 32'h00000000;
      queue_2_prd <= 6'h00;
      queue_2_psrc_0 <= 6'h00;
      queue_2_psrc_1 <= 6'h00;
      queue_2_imm <= 32'h00000000;
      queue_2_uop_muluOp <= MULUOp_mullo;
      queue_2_srcReady_0 <= 1'b0;
      queue_2_srcReady_1 <= 1'b0;
      queue_3_valid <= 1'b0;
      queue_3_robIdx <= 5'h00;
      queue_3_branchResult_targetPC <= 32'h00000000;
      queue_3_branchResult_branchResult <= 1'b0;
      queue_3_branchResult_predictFail <= 1'b0;
      queue_3_exceptionInfo_exception <= 1'b0;
      queue_3_exceptionInfo_eCode <= 6'h00;
      queue_3_exceptionInfo_eSubCode <= 1'b0;
      queue_3_pc <= 32'h00000000;
      queue_3_prd <= 6'h00;
      queue_3_psrc_0 <= 6'h00;
      queue_3_psrc_1 <= 6'h00;
      queue_3_imm <= 32'h00000000;
      queue_3_uop_muluOp <= MULUOp_mullo;
      queue_3_srcReady_0 <= 1'b0;
      queue_3_srcReady_1 <= 1'b0;
    end else begin
      queue_0_valid <= queueNext_0_valid;
      queue_0_robIdx <= queueNext_0_robIdx;
      queue_0_branchResult_targetPC <= queueNext_0_branchResult_targetPC;
      queue_0_branchResult_branchResult <= queueNext_0_branchResult_branchResult;
      queue_0_branchResult_predictFail <= queueNext_0_branchResult_predictFail;
      queue_0_exceptionInfo_exception <= queueNext_0_exceptionInfo_exception;
      queue_0_exceptionInfo_eCode <= queueNext_0_exceptionInfo_eCode;
      queue_0_exceptionInfo_eSubCode <= queueNext_0_exceptionInfo_eSubCode;
      queue_0_pc <= queueNext_0_pc;
      queue_0_prd <= queueNext_0_prd;
      queue_0_psrc_0 <= queueNext_0_psrc_0;
      queue_0_psrc_1 <= queueNext_0_psrc_1;
      queue_0_imm <= queueNext_0_imm;
      queue_0_uop_muluOp <= queueNext_0_uop_muluOp;
      queue_0_srcReady_0 <= queueNext_0_srcReady_0;
      queue_0_srcReady_1 <= queueNext_0_srcReady_1;
      queue_1_valid <= queueNext_1_valid;
      queue_1_robIdx <= queueNext_1_robIdx;
      queue_1_branchResult_targetPC <= queueNext_1_branchResult_targetPC;
      queue_1_branchResult_branchResult <= queueNext_1_branchResult_branchResult;
      queue_1_branchResult_predictFail <= queueNext_1_branchResult_predictFail;
      queue_1_exceptionInfo_exception <= queueNext_1_exceptionInfo_exception;
      queue_1_exceptionInfo_eCode <= queueNext_1_exceptionInfo_eCode;
      queue_1_exceptionInfo_eSubCode <= queueNext_1_exceptionInfo_eSubCode;
      queue_1_pc <= queueNext_1_pc;
      queue_1_prd <= queueNext_1_prd;
      queue_1_psrc_0 <= queueNext_1_psrc_0;
      queue_1_psrc_1 <= queueNext_1_psrc_1;
      queue_1_imm <= queueNext_1_imm;
      queue_1_uop_muluOp <= queueNext_1_uop_muluOp;
      queue_1_srcReady_0 <= queueNext_1_srcReady_0;
      queue_1_srcReady_1 <= queueNext_1_srcReady_1;
      queue_2_valid <= queueNext_2_valid;
      queue_2_robIdx <= queueNext_2_robIdx;
      queue_2_branchResult_targetPC <= queueNext_2_branchResult_targetPC;
      queue_2_branchResult_branchResult <= queueNext_2_branchResult_branchResult;
      queue_2_branchResult_predictFail <= queueNext_2_branchResult_predictFail;
      queue_2_exceptionInfo_exception <= queueNext_2_exceptionInfo_exception;
      queue_2_exceptionInfo_eCode <= queueNext_2_exceptionInfo_eCode;
      queue_2_exceptionInfo_eSubCode <= queueNext_2_exceptionInfo_eSubCode;
      queue_2_pc <= queueNext_2_pc;
      queue_2_prd <= queueNext_2_prd;
      queue_2_psrc_0 <= queueNext_2_psrc_0;
      queue_2_psrc_1 <= queueNext_2_psrc_1;
      queue_2_imm <= queueNext_2_imm;
      queue_2_uop_muluOp <= queueNext_2_uop_muluOp;
      queue_2_srcReady_0 <= queueNext_2_srcReady_0;
      queue_2_srcReady_1 <= queueNext_2_srcReady_1;
      queue_3_valid <= queueNext_3_valid;
      queue_3_robIdx <= queueNext_3_robIdx;
      queue_3_branchResult_targetPC <= queueNext_3_branchResult_targetPC;
      queue_3_branchResult_branchResult <= queueNext_3_branchResult_branchResult;
      queue_3_branchResult_predictFail <= queueNext_3_branchResult_predictFail;
      queue_3_exceptionInfo_exception <= queueNext_3_exceptionInfo_exception;
      queue_3_exceptionInfo_eCode <= queueNext_3_exceptionInfo_eCode;
      queue_3_exceptionInfo_eSubCode <= queueNext_3_exceptionInfo_eSubCode;
      queue_3_pc <= queueNext_3_pc;
      queue_3_prd <= queueNext_3_prd;
      queue_3_psrc_0 <= queueNext_3_psrc_0;
      queue_3_psrc_1 <= queueNext_3_psrc_1;
      queue_3_imm <= queueNext_3_imm;
      queue_3_uop_muluOp <= queueNext_3_uop_muluOp;
      queue_3_srcReady_0 <= queueNext_3_srcReady_0;
      queue_3_srcReady_1 <= queueNext_3_srcReady_1;
    end
  end


endmodule

module IssueQueue_1 (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [4:0]    io_input_payload_robIdx,
  input  wire [31:0]   io_input_payload_branchInfo_predictPC,
  input  wire          io_input_payload_branchInfo_predictResult,
  input  wire          io_input_payload_exceptionInfo_exception,
  input  wire [5:0]    io_input_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_input_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_payload_pc,
  input  wire [5:0]    io_input_payload_prd,
  input  wire [5:0]    io_input_payload_psrc_0,
  input  wire [5:0]    io_input_payload_psrc_1,
  input  wire [31:0]   io_input_payload_imm,
  input  wire [3:0]    io_input_payload_uop_aluOp,
  input  wire [1:0]    io_input_payload_uop_bruOp,
  input  wire [2:0]    io_input_payload_roop_aluROOp,
  input  wire [1:0]    io_input_payload_roop_cruROOp,
  input  wire          io_input_payload_srcReady_0,
  input  wire          io_input_payload_srcReady_1,
  output wire          io_csrInQueue,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [4:0]    io_output_payload_robIdx,
  output wire [31:0]   io_output_payload_branchInfo_predictPC,
  output wire          io_output_payload_branchInfo_predictResult,
  output wire          io_output_payload_exceptionInfo_exception,
  output wire [5:0]    io_output_payload_exceptionInfo_eCode,
  output wire [0:0]    io_output_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_output_payload_pc,
  output wire [5:0]    io_output_payload_prd,
  output wire [5:0]    io_output_payload_psrc_0,
  output wire [5:0]    io_output_payload_psrc_1,
  output wire [31:0]   io_output_payload_imm,
  output wire [3:0]    io_output_payload_uop_aluOp,
  output wire [1:0]    io_output_payload_uop_bruOp,
  output wire [2:0]    io_output_payload_roop_aluROOp,
  output wire [1:0]    io_output_payload_roop_cruROOp,
  input  wire [5:0]    io_writebackSignal_0,
  input  wire [5:0]    io_writebackSignal_1,
  input  wire [5:0]    io_writebackSignal_2,
  input  wire [5:0]    io_writebackSignal_3,
  input  wire [5:0]    io_writebackSignal_4,
  input  wire          io_earlyWakeup_0_valid,
  input  wire [5:0]    io_earlyWakeup_0_payload,
  input  wire          io_earlyWakeup_1_valid,
  input  wire [5:0]    io_earlyWakeup_1_payload,
  input  wire          io_earlyWakeup_2_valid,
  input  wire [5:0]    io_earlyWakeup_2_payload,
  input  wire          io_earlyWakeup_3_valid,
  input  wire [5:0]    io_earlyWakeup_3_payload,
  input  wire          io_earlyWakeup_4_valid,
  input  wire [5:0]    io_earlyWakeup_4_payload,
  input  wire          io_earlyWakeup_5_valid,
  input  wire [5:0]    io_earlyWakeup_5_payload,
  input  wire          io_earlyWakeup_6_valid,
  input  wire [5:0]    io_earlyWakeup_6_payload,
  input  wire          io_earlyWakeup_7_valid,
  input  wire [5:0]    io_earlyWakeup_7_payload,
  output wire          io_wakeOut_valid,
  output wire [5:0]    io_wakeOut_payload,
  input  wire          aclk,
  input  wire          cpuClockingArea_areaFlushReset_newReset
);
  localparam ALUOp_add = 4'd0;
  localparam ALUOp_sub = 4'd1;
  localparam ALUOp_slt = 4'd2;
  localparam ALUOp_sltu = 4'd3;
  localparam ALUOp_eq = 4'd4;
  localparam ALUOp_nor_1 = 4'd5;
  localparam ALUOp_and_1 = 4'd6;
  localparam ALUOp_or_1 = 4'd7;
  localparam ALUOp_xor_1 = 4'd8;
  localparam ALUOp_sll_1 = 4'd9;
  localparam ALUOp_srl_1 = 4'd10;
  localparam ALUOp_sra_1 = 4'd11;
  localparam ALUOp_passa = 4'd12;
  localparam ALUOp_passb = 4'd13;
  localparam BRUOp_nop = 2'd0;
  localparam BRUOp_add = 2'd1;
  localparam BRUOp_cadd = 2'd2;
  localparam BRUOp_ncadd = 2'd3;
  localparam ALUROOp_reg_1 = 3'd0;
  localparam ALUROOp_regimm = 3'd1;
  localparam ALUROOp_pcimm = 3'd2;
  localparam ALUROOp_csr = 3'd3;
  localparam ALUROOp_linkpc = 3'd4;
  localparam ALUROOp_linkreg = 3'd5;
  localparam CRUROOp_id = 2'd0;
  localparam CRUROOp_lo = 2'd1;
  localparam CRUROOp_hi = 2'd2;

  wire       [3:0]    _zz_readyToIssue_ohFirst_masked;
  wire       [4:0]    _zz_emptyEntry_ohFirst_masked;
  wire                _zz_appendEntry_srcReady_0;
  wire       [0:0]    _zz_appendEntry_srcReady_0_1;
  wire       [1:0]    _zz_appendEntry_srcReady_0_2;
  wire                _zz_appendEntry_srcReady_0_3;
  wire                _zz_appendEntry_srcReady_0_4;
  wire       [0:0]    _zz_appendEntry_srcReady_0_5;
  wire       [4:0]    _zz_appendEntry_srcReady_0_6;
  wire                _zz_appendEntry_srcReady_0_7;
  wire                _zz_appendEntry_srcReady_0_8;
  wire       [0:0]    _zz_appendEntry_srcReady_0_9;
  wire       [0:0]    _zz_appendEntry_srcReady_0_10;
  wire                _zz_appendEntry_srcReady_1;
  wire       [0:0]    _zz_appendEntry_srcReady_1_1;
  wire       [0:0]    _zz_appendEntry_srcReady_1_2;
  wire                _zz_appendEntry_srcReady_1_3;
  wire                _zz_appendEntry_srcReady_1_4;
  wire       [0:0]    _zz_appendEntry_srcReady_1_5;
  wire       [3:0]    _zz_appendEntry_srcReady_1_6;
  wire                _zz_updatedEntry_0_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_0_2;
  wire                _zz_updatedEntry_0_srcReady_0_3;
  wire                _zz_updatedEntry_0_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_0_5;
  wire       [3:0]    _zz_updatedEntry_0_srcReady_0_6;
  wire                _zz_updatedEntry_0_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_1_2;
  wire                _zz_updatedEntry_0_srcReady_1_3;
  wire                _zz_updatedEntry_0_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_1_5;
  wire       [3:0]    _zz_updatedEntry_0_srcReady_1_6;
  wire                _zz_updatedEntry_1_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_0_2;
  wire                _zz_updatedEntry_1_srcReady_0_3;
  wire                _zz_updatedEntry_1_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_0_5;
  wire       [3:0]    _zz_updatedEntry_1_srcReady_0_6;
  wire                _zz_updatedEntry_1_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_1_2;
  wire                _zz_updatedEntry_1_srcReady_1_3;
  wire                _zz_updatedEntry_1_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_1_5;
  wire       [3:0]    _zz_updatedEntry_1_srcReady_1_6;
  wire                _zz_updatedEntry_2_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_0_2;
  wire                _zz_updatedEntry_2_srcReady_0_3;
  wire                _zz_updatedEntry_2_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_0_5;
  wire       [3:0]    _zz_updatedEntry_2_srcReady_0_6;
  wire                _zz_updatedEntry_2_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_1_2;
  wire                _zz_updatedEntry_2_srcReady_1_3;
  wire                _zz_updatedEntry_2_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_1_5;
  wire       [3:0]    _zz_updatedEntry_2_srcReady_1_6;
  wire                _zz_updatedEntry_3_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_0_2;
  wire                _zz_updatedEntry_3_srcReady_0_3;
  wire                _zz_updatedEntry_3_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_0_5;
  wire       [3:0]    _zz_updatedEntry_3_srcReady_0_6;
  wire                _zz_updatedEntry_3_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_1_2;
  wire                _zz_updatedEntry_3_srcReady_1_3;
  wire                _zz_updatedEntry_3_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_1_5;
  wire       [3:0]    _zz_updatedEntry_3_srcReady_1_6;
  reg                 _zz_issueEntry_valid_4;
  reg        [4:0]    _zz_issueEntry_robIdx;
  reg        [31:0]   _zz_issueEntry_branchInfo_predictPC;
  reg                 _zz_issueEntry_branchInfo_predictResult;
  reg                 _zz_issueEntry_exceptionInfo_exception;
  reg        [5:0]    _zz_issueEntry_exceptionInfo_eCode;
  reg        [0:0]    _zz_issueEntry_exceptionInfo_eSubCode;
  reg        [31:0]   _zz_issueEntry_pc;
  reg        [5:0]    _zz_issueEntry_prd;
  reg        [5:0]    _zz_issueEntry_psrc_0;
  reg        [5:0]    _zz_issueEntry_psrc_1;
  reg        [31:0]   _zz_issueEntry_imm;
  reg        [3:0]    _zz_issueEntry_uop_aluOp;
  reg        [1:0]    _zz_issueEntry_uop_bruOp;
  reg        [2:0]    _zz_issueEntry_roop_aluROOp;
  reg        [1:0]    _zz_issueEntry_roop_cruROOp;
  reg                 _zz_issueEntry_srcReady_0;
  reg                 _zz_issueEntry_srcReady_1;
  reg                 queue_0_valid;
  reg        [4:0]    queue_0_robIdx;
  reg        [31:0]   queue_0_branchInfo_predictPC;
  reg                 queue_0_branchInfo_predictResult;
  reg                 queue_0_exceptionInfo_exception;
  reg        [5:0]    queue_0_exceptionInfo_eCode;
  reg        [0:0]    queue_0_exceptionInfo_eSubCode;
  reg        [31:0]   queue_0_pc;
  reg        [5:0]    queue_0_prd;
  reg        [5:0]    queue_0_psrc_0;
  reg        [5:0]    queue_0_psrc_1;
  reg        [31:0]   queue_0_imm;
  reg        [3:0]    queue_0_uop_aluOp;
  reg        [1:0]    queue_0_uop_bruOp;
  reg        [2:0]    queue_0_roop_aluROOp;
  reg        [1:0]    queue_0_roop_cruROOp;
  reg                 queue_0_srcReady_0;
  reg                 queue_0_srcReady_1;
  reg                 queue_1_valid;
  reg        [4:0]    queue_1_robIdx;
  reg        [31:0]   queue_1_branchInfo_predictPC;
  reg                 queue_1_branchInfo_predictResult;
  reg                 queue_1_exceptionInfo_exception;
  reg        [5:0]    queue_1_exceptionInfo_eCode;
  reg        [0:0]    queue_1_exceptionInfo_eSubCode;
  reg        [31:0]   queue_1_pc;
  reg        [5:0]    queue_1_prd;
  reg        [5:0]    queue_1_psrc_0;
  reg        [5:0]    queue_1_psrc_1;
  reg        [31:0]   queue_1_imm;
  reg        [3:0]    queue_1_uop_aluOp;
  reg        [1:0]    queue_1_uop_bruOp;
  reg        [2:0]    queue_1_roop_aluROOp;
  reg        [1:0]    queue_1_roop_cruROOp;
  reg                 queue_1_srcReady_0;
  reg                 queue_1_srcReady_1;
  reg                 queue_2_valid;
  reg        [4:0]    queue_2_robIdx;
  reg        [31:0]   queue_2_branchInfo_predictPC;
  reg                 queue_2_branchInfo_predictResult;
  reg                 queue_2_exceptionInfo_exception;
  reg        [5:0]    queue_2_exceptionInfo_eCode;
  reg        [0:0]    queue_2_exceptionInfo_eSubCode;
  reg        [31:0]   queue_2_pc;
  reg        [5:0]    queue_2_prd;
  reg        [5:0]    queue_2_psrc_0;
  reg        [5:0]    queue_2_psrc_1;
  reg        [31:0]   queue_2_imm;
  reg        [3:0]    queue_2_uop_aluOp;
  reg        [1:0]    queue_2_uop_bruOp;
  reg        [2:0]    queue_2_roop_aluROOp;
  reg        [1:0]    queue_2_roop_cruROOp;
  reg                 queue_2_srcReady_0;
  reg                 queue_2_srcReady_1;
  reg                 queue_3_valid;
  reg        [4:0]    queue_3_robIdx;
  reg        [31:0]   queue_3_branchInfo_predictPC;
  reg                 queue_3_branchInfo_predictResult;
  reg                 queue_3_exceptionInfo_exception;
  reg        [5:0]    queue_3_exceptionInfo_eCode;
  reg        [0:0]    queue_3_exceptionInfo_eSubCode;
  reg        [31:0]   queue_3_pc;
  reg        [5:0]    queue_3_prd;
  reg        [5:0]    queue_3_psrc_0;
  reg        [5:0]    queue_3_psrc_1;
  reg        [31:0]   queue_3_imm;
  reg        [3:0]    queue_3_uop_aluOp;
  reg        [1:0]    queue_3_uop_bruOp;
  reg        [2:0]    queue_3_roop_aluROOp;
  reg        [1:0]    queue_3_roop_cruROOp;
  reg                 queue_3_srcReady_0;
  reg                 queue_3_srcReady_1;
  reg        [3:0]    readyToIssue;
  wire       [3:0]    readyToIssue_ohFirst_input;
  wire       [3:0]    readyToIssue_ohFirst_masked;
  wire       [3:0]    issueVector;
  reg        [3:0]    shiftAhead;
  reg        [4:0]    emptyEntry;
  wire       [4:0]    emptyEntry_ohFirst_input;
  wire       [4:0]    emptyEntry_ohFirst_masked;
  wire       [4:0]    writeVector;
  wire                updatedEntry_0_valid;
  wire       [4:0]    updatedEntry_0_robIdx;
  wire       [31:0]   updatedEntry_0_branchInfo_predictPC;
  wire                updatedEntry_0_branchInfo_predictResult;
  wire                updatedEntry_0_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_0_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_0_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_0_pc;
  wire       [5:0]    updatedEntry_0_prd;
  wire       [5:0]    updatedEntry_0_psrc_0;
  wire       [5:0]    updatedEntry_0_psrc_1;
  wire       [31:0]   updatedEntry_0_imm;
  wire       [3:0]    updatedEntry_0_uop_aluOp;
  wire       [1:0]    updatedEntry_0_uop_bruOp;
  wire       [2:0]    updatedEntry_0_roop_aluROOp;
  wire       [1:0]    updatedEntry_0_roop_cruROOp;
  reg                 updatedEntry_0_srcReady_0;
  reg                 updatedEntry_0_srcReady_1;
  wire                updatedEntry_1_valid;
  wire       [4:0]    updatedEntry_1_robIdx;
  wire       [31:0]   updatedEntry_1_branchInfo_predictPC;
  wire                updatedEntry_1_branchInfo_predictResult;
  wire                updatedEntry_1_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_1_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_1_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_1_pc;
  wire       [5:0]    updatedEntry_1_prd;
  wire       [5:0]    updatedEntry_1_psrc_0;
  wire       [5:0]    updatedEntry_1_psrc_1;
  wire       [31:0]   updatedEntry_1_imm;
  wire       [3:0]    updatedEntry_1_uop_aluOp;
  wire       [1:0]    updatedEntry_1_uop_bruOp;
  wire       [2:0]    updatedEntry_1_roop_aluROOp;
  wire       [1:0]    updatedEntry_1_roop_cruROOp;
  reg                 updatedEntry_1_srcReady_0;
  reg                 updatedEntry_1_srcReady_1;
  wire                updatedEntry_2_valid;
  wire       [4:0]    updatedEntry_2_robIdx;
  wire       [31:0]   updatedEntry_2_branchInfo_predictPC;
  wire                updatedEntry_2_branchInfo_predictResult;
  wire                updatedEntry_2_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_2_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_2_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_2_pc;
  wire       [5:0]    updatedEntry_2_prd;
  wire       [5:0]    updatedEntry_2_psrc_0;
  wire       [5:0]    updatedEntry_2_psrc_1;
  wire       [31:0]   updatedEntry_2_imm;
  wire       [3:0]    updatedEntry_2_uop_aluOp;
  wire       [1:0]    updatedEntry_2_uop_bruOp;
  wire       [2:0]    updatedEntry_2_roop_aluROOp;
  wire       [1:0]    updatedEntry_2_roop_cruROOp;
  reg                 updatedEntry_2_srcReady_0;
  reg                 updatedEntry_2_srcReady_1;
  wire                updatedEntry_3_valid;
  wire       [4:0]    updatedEntry_3_robIdx;
  wire       [31:0]   updatedEntry_3_branchInfo_predictPC;
  wire                updatedEntry_3_branchInfo_predictResult;
  wire                updatedEntry_3_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_3_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_3_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_3_pc;
  wire       [5:0]    updatedEntry_3_prd;
  wire       [5:0]    updatedEntry_3_psrc_0;
  wire       [5:0]    updatedEntry_3_psrc_1;
  wire       [31:0]   updatedEntry_3_imm;
  wire       [3:0]    updatedEntry_3_uop_aluOp;
  wire       [1:0]    updatedEntry_3_uop_bruOp;
  wire       [2:0]    updatedEntry_3_roop_aluROOp;
  wire       [1:0]    updatedEntry_3_roop_cruROOp;
  reg                 updatedEntry_3_srcReady_0;
  reg                 updatedEntry_3_srcReady_1;
  wire                appendEntry_valid;
  wire       [4:0]    appendEntry_robIdx;
  wire       [31:0]   appendEntry_branchInfo_predictPC;
  wire                appendEntry_branchInfo_predictResult;
  wire                appendEntry_exceptionInfo_exception;
  wire       [5:0]    appendEntry_exceptionInfo_eCode;
  wire       [0:0]    appendEntry_exceptionInfo_eSubCode;
  wire       [31:0]   appendEntry_pc;
  wire       [5:0]    appendEntry_prd;
  wire       [5:0]    appendEntry_psrc_0;
  wire       [5:0]    appendEntry_psrc_1;
  wire       [31:0]   appendEntry_imm;
  wire       [3:0]    appendEntry_uop_aluOp;
  wire       [1:0]    appendEntry_uop_bruOp;
  wire       [2:0]    appendEntry_roop_aluROOp;
  wire       [1:0]    appendEntry_roop_cruROOp;
  wire                appendEntry_srcReady_0;
  wire                appendEntry_srcReady_1;
  reg                 queueNext_0_valid;
  reg        [4:0]    queueNext_0_robIdx;
  reg        [31:0]   queueNext_0_branchInfo_predictPC;
  reg                 queueNext_0_branchInfo_predictResult;
  reg                 queueNext_0_exceptionInfo_exception;
  reg        [5:0]    queueNext_0_exceptionInfo_eCode;
  reg        [0:0]    queueNext_0_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_0_pc;
  reg        [5:0]    queueNext_0_prd;
  reg        [5:0]    queueNext_0_psrc_0;
  reg        [5:0]    queueNext_0_psrc_1;
  reg        [31:0]   queueNext_0_imm;
  reg        [3:0]    queueNext_0_uop_aluOp;
  reg        [1:0]    queueNext_0_uop_bruOp;
  reg        [2:0]    queueNext_0_roop_aluROOp;
  reg        [1:0]    queueNext_0_roop_cruROOp;
  reg                 queueNext_0_srcReady_0;
  reg                 queueNext_0_srcReady_1;
  reg                 queueNext_1_valid;
  reg        [4:0]    queueNext_1_robIdx;
  reg        [31:0]   queueNext_1_branchInfo_predictPC;
  reg                 queueNext_1_branchInfo_predictResult;
  reg                 queueNext_1_exceptionInfo_exception;
  reg        [5:0]    queueNext_1_exceptionInfo_eCode;
  reg        [0:0]    queueNext_1_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_1_pc;
  reg        [5:0]    queueNext_1_prd;
  reg        [5:0]    queueNext_1_psrc_0;
  reg        [5:0]    queueNext_1_psrc_1;
  reg        [31:0]   queueNext_1_imm;
  reg        [3:0]    queueNext_1_uop_aluOp;
  reg        [1:0]    queueNext_1_uop_bruOp;
  reg        [2:0]    queueNext_1_roop_aluROOp;
  reg        [1:0]    queueNext_1_roop_cruROOp;
  reg                 queueNext_1_srcReady_0;
  reg                 queueNext_1_srcReady_1;
  reg                 queueNext_2_valid;
  reg        [4:0]    queueNext_2_robIdx;
  reg        [31:0]   queueNext_2_branchInfo_predictPC;
  reg                 queueNext_2_branchInfo_predictResult;
  reg                 queueNext_2_exceptionInfo_exception;
  reg        [5:0]    queueNext_2_exceptionInfo_eCode;
  reg        [0:0]    queueNext_2_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_2_pc;
  reg        [5:0]    queueNext_2_prd;
  reg        [5:0]    queueNext_2_psrc_0;
  reg        [5:0]    queueNext_2_psrc_1;
  reg        [31:0]   queueNext_2_imm;
  reg        [3:0]    queueNext_2_uop_aluOp;
  reg        [1:0]    queueNext_2_uop_bruOp;
  reg        [2:0]    queueNext_2_roop_aluROOp;
  reg        [1:0]    queueNext_2_roop_cruROOp;
  reg                 queueNext_2_srcReady_0;
  reg                 queueNext_2_srcReady_1;
  reg                 queueNext_3_valid;
  reg        [4:0]    queueNext_3_robIdx;
  reg        [31:0]   queueNext_3_branchInfo_predictPC;
  reg                 queueNext_3_branchInfo_predictResult;
  reg                 queueNext_3_exceptionInfo_exception;
  reg        [5:0]    queueNext_3_exceptionInfo_eCode;
  reg        [0:0]    queueNext_3_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_3_pc;
  reg        [5:0]    queueNext_3_prd;
  reg        [5:0]    queueNext_3_psrc_0;
  reg        [5:0]    queueNext_3_psrc_1;
  reg        [31:0]   queueNext_3_imm;
  reg        [3:0]    queueNext_3_uop_aluOp;
  reg        [1:0]    queueNext_3_uop_bruOp;
  reg        [2:0]    queueNext_3_roop_aluROOp;
  reg        [1:0]    queueNext_3_roop_cruROOp;
  reg                 queueNext_3_srcReady_0;
  reg                 queueNext_3_srcReady_1;
  wire                when_IssueQueue_l81;
  wire                when_IssueQueue_l83;
  wire                when_IssueQueue_l96;
  wire                when_IssueQueue_l81_1;
  wire                when_IssueQueue_l83_1;
  wire                when_IssueQueue_l96_1;
  wire                when_IssueQueue_l81_2;
  wire                when_IssueQueue_l83_2;
  wire                when_IssueQueue_l96_2;
  wire                when_IssueQueue_l81_3;
  wire                when_IssueQueue_l89;
  wire                when_IssueQueue_l96_3;
  reg        [3:0]    _zz_io_csrInQueue;
  wire                io_output_fire;
  wire                _zz_issueEntry_valid;
  wire                _zz_issueEntry_valid_1;
  wire                _zz_issueEntry_valid_2;
  wire       [1:0]    _zz_issueEntry_valid_3;
  wire                issueEntry_valid;
  wire       [4:0]    issueEntry_robIdx;
  wire       [31:0]   issueEntry_branchInfo_predictPC;
  wire                issueEntry_branchInfo_predictResult;
  wire                issueEntry_exceptionInfo_exception;
  wire       [5:0]    issueEntry_exceptionInfo_eCode;
  wire       [0:0]    issueEntry_exceptionInfo_eSubCode;
  wire       [31:0]   issueEntry_pc;
  wire       [5:0]    issueEntry_prd;
  wire       [5:0]    issueEntry_psrc_0;
  wire       [5:0]    issueEntry_psrc_1;
  wire       [31:0]   issueEntry_imm;
  wire       [3:0]    issueEntry_uop_aluOp;
  wire       [1:0]    issueEntry_uop_bruOp;
  wire       [2:0]    issueEntry_roop_aluROOp;
  wire       [1:0]    issueEntry_roop_cruROOp;
  wire                issueEntry_srcReady_0;
  wire                issueEntry_srcReady_1;
  `ifndef SYNTHESIS
  reg [39:0] io_input_payload_uop_aluOp_string;
  reg [39:0] io_input_payload_uop_bruOp_string;
  reg [55:0] io_input_payload_roop_aluROOp_string;
  reg [15:0] io_input_payload_roop_cruROOp_string;
  reg [39:0] io_output_payload_uop_aluOp_string;
  reg [39:0] io_output_payload_uop_bruOp_string;
  reg [55:0] io_output_payload_roop_aluROOp_string;
  reg [15:0] io_output_payload_roop_cruROOp_string;
  reg [39:0] queue_0_uop_aluOp_string;
  reg [39:0] queue_0_uop_bruOp_string;
  reg [55:0] queue_0_roop_aluROOp_string;
  reg [15:0] queue_0_roop_cruROOp_string;
  reg [39:0] queue_1_uop_aluOp_string;
  reg [39:0] queue_1_uop_bruOp_string;
  reg [55:0] queue_1_roop_aluROOp_string;
  reg [15:0] queue_1_roop_cruROOp_string;
  reg [39:0] queue_2_uop_aluOp_string;
  reg [39:0] queue_2_uop_bruOp_string;
  reg [55:0] queue_2_roop_aluROOp_string;
  reg [15:0] queue_2_roop_cruROOp_string;
  reg [39:0] queue_3_uop_aluOp_string;
  reg [39:0] queue_3_uop_bruOp_string;
  reg [55:0] queue_3_roop_aluROOp_string;
  reg [15:0] queue_3_roop_cruROOp_string;
  reg [39:0] updatedEntry_0_uop_aluOp_string;
  reg [39:0] updatedEntry_0_uop_bruOp_string;
  reg [55:0] updatedEntry_0_roop_aluROOp_string;
  reg [15:0] updatedEntry_0_roop_cruROOp_string;
  reg [39:0] updatedEntry_1_uop_aluOp_string;
  reg [39:0] updatedEntry_1_uop_bruOp_string;
  reg [55:0] updatedEntry_1_roop_aluROOp_string;
  reg [15:0] updatedEntry_1_roop_cruROOp_string;
  reg [39:0] updatedEntry_2_uop_aluOp_string;
  reg [39:0] updatedEntry_2_uop_bruOp_string;
  reg [55:0] updatedEntry_2_roop_aluROOp_string;
  reg [15:0] updatedEntry_2_roop_cruROOp_string;
  reg [39:0] updatedEntry_3_uop_aluOp_string;
  reg [39:0] updatedEntry_3_uop_bruOp_string;
  reg [55:0] updatedEntry_3_roop_aluROOp_string;
  reg [15:0] updatedEntry_3_roop_cruROOp_string;
  reg [39:0] appendEntry_uop_aluOp_string;
  reg [39:0] appendEntry_uop_bruOp_string;
  reg [55:0] appendEntry_roop_aluROOp_string;
  reg [15:0] appendEntry_roop_cruROOp_string;
  reg [39:0] queueNext_0_uop_aluOp_string;
  reg [39:0] queueNext_0_uop_bruOp_string;
  reg [55:0] queueNext_0_roop_aluROOp_string;
  reg [15:0] queueNext_0_roop_cruROOp_string;
  reg [39:0] queueNext_1_uop_aluOp_string;
  reg [39:0] queueNext_1_uop_bruOp_string;
  reg [55:0] queueNext_1_roop_aluROOp_string;
  reg [15:0] queueNext_1_roop_cruROOp_string;
  reg [39:0] queueNext_2_uop_aluOp_string;
  reg [39:0] queueNext_2_uop_bruOp_string;
  reg [55:0] queueNext_2_roop_aluROOp_string;
  reg [15:0] queueNext_2_roop_cruROOp_string;
  reg [39:0] queueNext_3_uop_aluOp_string;
  reg [39:0] queueNext_3_uop_bruOp_string;
  reg [55:0] queueNext_3_roop_aluROOp_string;
  reg [15:0] queueNext_3_roop_cruROOp_string;
  reg [39:0] issueEntry_uop_aluOp_string;
  reg [39:0] issueEntry_uop_bruOp_string;
  reg [55:0] issueEntry_roop_aluROOp_string;
  reg [15:0] issueEntry_roop_cruROOp_string;
  `endif


  assign _zz_readyToIssue_ohFirst_masked = (readyToIssue_ohFirst_input - 4'b0001);
  assign _zz_emptyEntry_ohFirst_masked = (emptyEntry_ohFirst_input - 5'h01);
  assign _zz_appendEntry_srcReady_0 = (io_input_payload_psrc_0 == io_writebackSignal_3);
  assign _zz_appendEntry_srcReady_0_1 = (io_input_payload_psrc_0 == io_writebackSignal_2);
  assign _zz_appendEntry_srcReady_0_2 = {(io_input_payload_psrc_0 == io_writebackSignal_1),(io_input_payload_psrc_0 == io_writebackSignal_0)};
  assign _zz_appendEntry_srcReady_0_3 = (io_input_payload_psrc_0 == io_earlyWakeup_7_payload);
  assign _zz_appendEntry_srcReady_0_4 = ((io_input_payload_psrc_0 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid);
  assign _zz_appendEntry_srcReady_0_5 = ((io_input_payload_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_appendEntry_srcReady_0_6 = {((io_input_payload_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid),{(_zz_appendEntry_srcReady_0_7 && io_earlyWakeup_3_valid),{_zz_appendEntry_srcReady_0_8,{_zz_appendEntry_srcReady_0_9,_zz_appendEntry_srcReady_0_10}}}};
  assign _zz_appendEntry_srcReady_0_7 = (io_input_payload_psrc_0 == io_earlyWakeup_3_payload);
  assign _zz_appendEntry_srcReady_0_8 = ((io_input_payload_psrc_0 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid);
  assign _zz_appendEntry_srcReady_0_9 = ((io_input_payload_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid);
  assign _zz_appendEntry_srcReady_0_10 = ((io_input_payload_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid);
  assign _zz_appendEntry_srcReady_1 = (io_input_payload_psrc_1 == io_writebackSignal_2);
  assign _zz_appendEntry_srcReady_1_1 = (io_input_payload_psrc_1 == io_writebackSignal_1);
  assign _zz_appendEntry_srcReady_1_2 = (io_input_payload_psrc_1 == io_writebackSignal_0);
  assign _zz_appendEntry_srcReady_1_3 = (io_input_payload_psrc_1 == io_earlyWakeup_6_payload);
  assign _zz_appendEntry_srcReady_1_4 = ((io_input_payload_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_appendEntry_srcReady_1_5 = ((io_input_payload_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_appendEntry_srcReady_1_6 = {((io_input_payload_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((io_input_payload_psrc_1 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((io_input_payload_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((io_input_payload_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_0_srcReady_0 = (queue_0_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_0_srcReady_0_1 = (queue_0_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_0_srcReady_0_2 = (queue_0_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_0_srcReady_0_3 = (queue_0_psrc_0 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_0_srcReady_0_4 = ((queue_0_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_0_srcReady_0_5 = ((queue_0_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_0_srcReady_0_6 = {((queue_0_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_0_psrc_0 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_0_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_0_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_0_srcReady_1 = (queue_0_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_0_srcReady_1_1 = (queue_0_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_0_srcReady_1_2 = (queue_0_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_0_srcReady_1_3 = (queue_0_psrc_1 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_0_srcReady_1_4 = ((queue_0_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_0_srcReady_1_5 = ((queue_0_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_0_srcReady_1_6 = {((queue_0_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_0_psrc_1 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_0_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_0_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_1_srcReady_0 = (queue_1_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_1_srcReady_0_1 = (queue_1_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_1_srcReady_0_2 = (queue_1_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_1_srcReady_0_3 = (queue_1_psrc_0 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_1_srcReady_0_4 = ((queue_1_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_1_srcReady_0_5 = ((queue_1_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_1_srcReady_0_6 = {((queue_1_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_1_psrc_0 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_1_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_1_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_1_srcReady_1 = (queue_1_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_1_srcReady_1_1 = (queue_1_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_1_srcReady_1_2 = (queue_1_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_1_srcReady_1_3 = (queue_1_psrc_1 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_1_srcReady_1_4 = ((queue_1_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_1_srcReady_1_5 = ((queue_1_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_1_srcReady_1_6 = {((queue_1_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_1_psrc_1 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_1_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_1_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_2_srcReady_0 = (queue_2_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_2_srcReady_0_1 = (queue_2_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_2_srcReady_0_2 = (queue_2_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_2_srcReady_0_3 = (queue_2_psrc_0 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_2_srcReady_0_4 = ((queue_2_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_2_srcReady_0_5 = ((queue_2_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_2_srcReady_0_6 = {((queue_2_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_2_psrc_0 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_2_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_2_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_2_srcReady_1 = (queue_2_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_2_srcReady_1_1 = (queue_2_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_2_srcReady_1_2 = (queue_2_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_2_srcReady_1_3 = (queue_2_psrc_1 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_2_srcReady_1_4 = ((queue_2_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_2_srcReady_1_5 = ((queue_2_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_2_srcReady_1_6 = {((queue_2_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_2_psrc_1 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_2_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_2_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_3_srcReady_0 = (queue_3_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_3_srcReady_0_1 = (queue_3_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_3_srcReady_0_2 = (queue_3_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_3_srcReady_0_3 = (queue_3_psrc_0 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_3_srcReady_0_4 = ((queue_3_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_3_srcReady_0_5 = ((queue_3_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_3_srcReady_0_6 = {((queue_3_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_3_psrc_0 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_3_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_3_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_3_srcReady_1 = (queue_3_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_3_srcReady_1_1 = (queue_3_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_3_srcReady_1_2 = (queue_3_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_3_srcReady_1_3 = (queue_3_psrc_1 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_3_srcReady_1_4 = ((queue_3_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_3_srcReady_1_5 = ((queue_3_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_3_srcReady_1_6 = {((queue_3_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_3_psrc_1 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_3_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_3_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  always @(*) begin
    case(_zz_issueEntry_valid_3)
      2'b00 : begin
        _zz_issueEntry_valid_4 = queue_0_valid;
        _zz_issueEntry_robIdx = queue_0_robIdx;
        _zz_issueEntry_branchInfo_predictPC = queue_0_branchInfo_predictPC;
        _zz_issueEntry_branchInfo_predictResult = queue_0_branchInfo_predictResult;
        _zz_issueEntry_exceptionInfo_exception = queue_0_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_0_pc;
        _zz_issueEntry_prd = queue_0_prd;
        _zz_issueEntry_psrc_0 = queue_0_psrc_0;
        _zz_issueEntry_psrc_1 = queue_0_psrc_1;
        _zz_issueEntry_imm = queue_0_imm;
        _zz_issueEntry_uop_aluOp = queue_0_uop_aluOp;
        _zz_issueEntry_uop_bruOp = queue_0_uop_bruOp;
        _zz_issueEntry_roop_aluROOp = queue_0_roop_aluROOp;
        _zz_issueEntry_roop_cruROOp = queue_0_roop_cruROOp;
        _zz_issueEntry_srcReady_0 = queue_0_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_0_srcReady_1;
      end
      2'b01 : begin
        _zz_issueEntry_valid_4 = queue_1_valid;
        _zz_issueEntry_robIdx = queue_1_robIdx;
        _zz_issueEntry_branchInfo_predictPC = queue_1_branchInfo_predictPC;
        _zz_issueEntry_branchInfo_predictResult = queue_1_branchInfo_predictResult;
        _zz_issueEntry_exceptionInfo_exception = queue_1_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_1_pc;
        _zz_issueEntry_prd = queue_1_prd;
        _zz_issueEntry_psrc_0 = queue_1_psrc_0;
        _zz_issueEntry_psrc_1 = queue_1_psrc_1;
        _zz_issueEntry_imm = queue_1_imm;
        _zz_issueEntry_uop_aluOp = queue_1_uop_aluOp;
        _zz_issueEntry_uop_bruOp = queue_1_uop_bruOp;
        _zz_issueEntry_roop_aluROOp = queue_1_roop_aluROOp;
        _zz_issueEntry_roop_cruROOp = queue_1_roop_cruROOp;
        _zz_issueEntry_srcReady_0 = queue_1_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_1_srcReady_1;
      end
      2'b10 : begin
        _zz_issueEntry_valid_4 = queue_2_valid;
        _zz_issueEntry_robIdx = queue_2_robIdx;
        _zz_issueEntry_branchInfo_predictPC = queue_2_branchInfo_predictPC;
        _zz_issueEntry_branchInfo_predictResult = queue_2_branchInfo_predictResult;
        _zz_issueEntry_exceptionInfo_exception = queue_2_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_2_pc;
        _zz_issueEntry_prd = queue_2_prd;
        _zz_issueEntry_psrc_0 = queue_2_psrc_0;
        _zz_issueEntry_psrc_1 = queue_2_psrc_1;
        _zz_issueEntry_imm = queue_2_imm;
        _zz_issueEntry_uop_aluOp = queue_2_uop_aluOp;
        _zz_issueEntry_uop_bruOp = queue_2_uop_bruOp;
        _zz_issueEntry_roop_aluROOp = queue_2_roop_aluROOp;
        _zz_issueEntry_roop_cruROOp = queue_2_roop_cruROOp;
        _zz_issueEntry_srcReady_0 = queue_2_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_2_srcReady_1;
      end
      default : begin
        _zz_issueEntry_valid_4 = queue_3_valid;
        _zz_issueEntry_robIdx = queue_3_robIdx;
        _zz_issueEntry_branchInfo_predictPC = queue_3_branchInfo_predictPC;
        _zz_issueEntry_branchInfo_predictResult = queue_3_branchInfo_predictResult;
        _zz_issueEntry_exceptionInfo_exception = queue_3_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_3_pc;
        _zz_issueEntry_prd = queue_3_prd;
        _zz_issueEntry_psrc_0 = queue_3_psrc_0;
        _zz_issueEntry_psrc_1 = queue_3_psrc_1;
        _zz_issueEntry_imm = queue_3_imm;
        _zz_issueEntry_uop_aluOp = queue_3_uop_aluOp;
        _zz_issueEntry_uop_bruOp = queue_3_uop_bruOp;
        _zz_issueEntry_roop_aluROOp = queue_3_roop_aluROOp;
        _zz_issueEntry_roop_cruROOp = queue_3_roop_cruROOp;
        _zz_issueEntry_srcReady_0 = queue_3_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_3_srcReady_1;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_uop_aluOp)
      ALUOp_add : io_input_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_input_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_input_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_input_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_input_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_input_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_input_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_input_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_input_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_input_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_input_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_input_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_input_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_input_payload_uop_aluOp_string = "passb";
      default : io_input_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_input_payload_uop_bruOp)
      BRUOp_nop : io_input_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_input_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_input_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_input_payload_uop_bruOp_string = "ncadd";
      default : io_input_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_input_payload_roop_aluROOp)
      ALUROOp_reg_1 : io_input_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : io_input_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : io_input_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : io_input_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : io_input_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : io_input_payload_roop_aluROOp_string = "linkreg";
      default : io_input_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_input_payload_roop_cruROOp)
      CRUROOp_id : io_input_payload_roop_cruROOp_string = "id";
      CRUROOp_lo : io_input_payload_roop_cruROOp_string = "lo";
      CRUROOp_hi : io_input_payload_roop_cruROOp_string = "hi";
      default : io_input_payload_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(io_output_payload_uop_aluOp)
      ALUOp_add : io_output_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_output_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_output_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_output_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_output_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_output_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_output_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_output_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_output_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_output_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_output_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_output_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_output_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_output_payload_uop_aluOp_string = "passb";
      default : io_output_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_uop_bruOp)
      BRUOp_nop : io_output_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_output_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_output_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_output_payload_uop_bruOp_string = "ncadd";
      default : io_output_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_roop_aluROOp)
      ALUROOp_reg_1 : io_output_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : io_output_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : io_output_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : io_output_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : io_output_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : io_output_payload_roop_aluROOp_string = "linkreg";
      default : io_output_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_roop_cruROOp)
      CRUROOp_id : io_output_payload_roop_cruROOp_string = "id";
      CRUROOp_lo : io_output_payload_roop_cruROOp_string = "lo";
      CRUROOp_hi : io_output_payload_roop_cruROOp_string = "hi";
      default : io_output_payload_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(queue_0_uop_aluOp)
      ALUOp_add : queue_0_uop_aluOp_string = "add  ";
      ALUOp_sub : queue_0_uop_aluOp_string = "sub  ";
      ALUOp_slt : queue_0_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queue_0_uop_aluOp_string = "sltu ";
      ALUOp_eq : queue_0_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queue_0_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queue_0_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queue_0_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queue_0_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queue_0_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queue_0_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queue_0_uop_aluOp_string = "sra_1";
      ALUOp_passa : queue_0_uop_aluOp_string = "passa";
      ALUOp_passb : queue_0_uop_aluOp_string = "passb";
      default : queue_0_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_0_uop_bruOp)
      BRUOp_nop : queue_0_uop_bruOp_string = "nop  ";
      BRUOp_add : queue_0_uop_bruOp_string = "add  ";
      BRUOp_cadd : queue_0_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queue_0_uop_bruOp_string = "ncadd";
      default : queue_0_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_0_roop_aluROOp)
      ALUROOp_reg_1 : queue_0_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queue_0_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queue_0_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queue_0_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queue_0_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queue_0_roop_aluROOp_string = "linkreg";
      default : queue_0_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_0_roop_cruROOp)
      CRUROOp_id : queue_0_roop_cruROOp_string = "id";
      CRUROOp_lo : queue_0_roop_cruROOp_string = "lo";
      CRUROOp_hi : queue_0_roop_cruROOp_string = "hi";
      default : queue_0_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(queue_1_uop_aluOp)
      ALUOp_add : queue_1_uop_aluOp_string = "add  ";
      ALUOp_sub : queue_1_uop_aluOp_string = "sub  ";
      ALUOp_slt : queue_1_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queue_1_uop_aluOp_string = "sltu ";
      ALUOp_eq : queue_1_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queue_1_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queue_1_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queue_1_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queue_1_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queue_1_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queue_1_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queue_1_uop_aluOp_string = "sra_1";
      ALUOp_passa : queue_1_uop_aluOp_string = "passa";
      ALUOp_passb : queue_1_uop_aluOp_string = "passb";
      default : queue_1_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_1_uop_bruOp)
      BRUOp_nop : queue_1_uop_bruOp_string = "nop  ";
      BRUOp_add : queue_1_uop_bruOp_string = "add  ";
      BRUOp_cadd : queue_1_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queue_1_uop_bruOp_string = "ncadd";
      default : queue_1_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_1_roop_aluROOp)
      ALUROOp_reg_1 : queue_1_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queue_1_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queue_1_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queue_1_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queue_1_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queue_1_roop_aluROOp_string = "linkreg";
      default : queue_1_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_1_roop_cruROOp)
      CRUROOp_id : queue_1_roop_cruROOp_string = "id";
      CRUROOp_lo : queue_1_roop_cruROOp_string = "lo";
      CRUROOp_hi : queue_1_roop_cruROOp_string = "hi";
      default : queue_1_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(queue_2_uop_aluOp)
      ALUOp_add : queue_2_uop_aluOp_string = "add  ";
      ALUOp_sub : queue_2_uop_aluOp_string = "sub  ";
      ALUOp_slt : queue_2_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queue_2_uop_aluOp_string = "sltu ";
      ALUOp_eq : queue_2_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queue_2_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queue_2_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queue_2_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queue_2_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queue_2_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queue_2_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queue_2_uop_aluOp_string = "sra_1";
      ALUOp_passa : queue_2_uop_aluOp_string = "passa";
      ALUOp_passb : queue_2_uop_aluOp_string = "passb";
      default : queue_2_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_2_uop_bruOp)
      BRUOp_nop : queue_2_uop_bruOp_string = "nop  ";
      BRUOp_add : queue_2_uop_bruOp_string = "add  ";
      BRUOp_cadd : queue_2_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queue_2_uop_bruOp_string = "ncadd";
      default : queue_2_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_2_roop_aluROOp)
      ALUROOp_reg_1 : queue_2_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queue_2_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queue_2_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queue_2_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queue_2_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queue_2_roop_aluROOp_string = "linkreg";
      default : queue_2_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_2_roop_cruROOp)
      CRUROOp_id : queue_2_roop_cruROOp_string = "id";
      CRUROOp_lo : queue_2_roop_cruROOp_string = "lo";
      CRUROOp_hi : queue_2_roop_cruROOp_string = "hi";
      default : queue_2_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(queue_3_uop_aluOp)
      ALUOp_add : queue_3_uop_aluOp_string = "add  ";
      ALUOp_sub : queue_3_uop_aluOp_string = "sub  ";
      ALUOp_slt : queue_3_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queue_3_uop_aluOp_string = "sltu ";
      ALUOp_eq : queue_3_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queue_3_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queue_3_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queue_3_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queue_3_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queue_3_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queue_3_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queue_3_uop_aluOp_string = "sra_1";
      ALUOp_passa : queue_3_uop_aluOp_string = "passa";
      ALUOp_passb : queue_3_uop_aluOp_string = "passb";
      default : queue_3_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_3_uop_bruOp)
      BRUOp_nop : queue_3_uop_bruOp_string = "nop  ";
      BRUOp_add : queue_3_uop_bruOp_string = "add  ";
      BRUOp_cadd : queue_3_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queue_3_uop_bruOp_string = "ncadd";
      default : queue_3_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_3_roop_aluROOp)
      ALUROOp_reg_1 : queue_3_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queue_3_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queue_3_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queue_3_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queue_3_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queue_3_roop_aluROOp_string = "linkreg";
      default : queue_3_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_3_roop_cruROOp)
      CRUROOp_id : queue_3_roop_cruROOp_string = "id";
      CRUROOp_lo : queue_3_roop_cruROOp_string = "lo";
      CRUROOp_hi : queue_3_roop_cruROOp_string = "hi";
      default : queue_3_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_uop_aluOp)
      ALUOp_add : updatedEntry_0_uop_aluOp_string = "add  ";
      ALUOp_sub : updatedEntry_0_uop_aluOp_string = "sub  ";
      ALUOp_slt : updatedEntry_0_uop_aluOp_string = "slt  ";
      ALUOp_sltu : updatedEntry_0_uop_aluOp_string = "sltu ";
      ALUOp_eq : updatedEntry_0_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : updatedEntry_0_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : updatedEntry_0_uop_aluOp_string = "and_1";
      ALUOp_or_1 : updatedEntry_0_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : updatedEntry_0_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : updatedEntry_0_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : updatedEntry_0_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : updatedEntry_0_uop_aluOp_string = "sra_1";
      ALUOp_passa : updatedEntry_0_uop_aluOp_string = "passa";
      ALUOp_passb : updatedEntry_0_uop_aluOp_string = "passb";
      default : updatedEntry_0_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_uop_bruOp)
      BRUOp_nop : updatedEntry_0_uop_bruOp_string = "nop  ";
      BRUOp_add : updatedEntry_0_uop_bruOp_string = "add  ";
      BRUOp_cadd : updatedEntry_0_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : updatedEntry_0_uop_bruOp_string = "ncadd";
      default : updatedEntry_0_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_roop_aluROOp)
      ALUROOp_reg_1 : updatedEntry_0_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : updatedEntry_0_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : updatedEntry_0_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : updatedEntry_0_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : updatedEntry_0_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : updatedEntry_0_roop_aluROOp_string = "linkreg";
      default : updatedEntry_0_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_roop_cruROOp)
      CRUROOp_id : updatedEntry_0_roop_cruROOp_string = "id";
      CRUROOp_lo : updatedEntry_0_roop_cruROOp_string = "lo";
      CRUROOp_hi : updatedEntry_0_roop_cruROOp_string = "hi";
      default : updatedEntry_0_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_uop_aluOp)
      ALUOp_add : updatedEntry_1_uop_aluOp_string = "add  ";
      ALUOp_sub : updatedEntry_1_uop_aluOp_string = "sub  ";
      ALUOp_slt : updatedEntry_1_uop_aluOp_string = "slt  ";
      ALUOp_sltu : updatedEntry_1_uop_aluOp_string = "sltu ";
      ALUOp_eq : updatedEntry_1_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : updatedEntry_1_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : updatedEntry_1_uop_aluOp_string = "and_1";
      ALUOp_or_1 : updatedEntry_1_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : updatedEntry_1_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : updatedEntry_1_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : updatedEntry_1_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : updatedEntry_1_uop_aluOp_string = "sra_1";
      ALUOp_passa : updatedEntry_1_uop_aluOp_string = "passa";
      ALUOp_passb : updatedEntry_1_uop_aluOp_string = "passb";
      default : updatedEntry_1_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_uop_bruOp)
      BRUOp_nop : updatedEntry_1_uop_bruOp_string = "nop  ";
      BRUOp_add : updatedEntry_1_uop_bruOp_string = "add  ";
      BRUOp_cadd : updatedEntry_1_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : updatedEntry_1_uop_bruOp_string = "ncadd";
      default : updatedEntry_1_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_roop_aluROOp)
      ALUROOp_reg_1 : updatedEntry_1_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : updatedEntry_1_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : updatedEntry_1_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : updatedEntry_1_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : updatedEntry_1_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : updatedEntry_1_roop_aluROOp_string = "linkreg";
      default : updatedEntry_1_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_roop_cruROOp)
      CRUROOp_id : updatedEntry_1_roop_cruROOp_string = "id";
      CRUROOp_lo : updatedEntry_1_roop_cruROOp_string = "lo";
      CRUROOp_hi : updatedEntry_1_roop_cruROOp_string = "hi";
      default : updatedEntry_1_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_uop_aluOp)
      ALUOp_add : updatedEntry_2_uop_aluOp_string = "add  ";
      ALUOp_sub : updatedEntry_2_uop_aluOp_string = "sub  ";
      ALUOp_slt : updatedEntry_2_uop_aluOp_string = "slt  ";
      ALUOp_sltu : updatedEntry_2_uop_aluOp_string = "sltu ";
      ALUOp_eq : updatedEntry_2_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : updatedEntry_2_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : updatedEntry_2_uop_aluOp_string = "and_1";
      ALUOp_or_1 : updatedEntry_2_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : updatedEntry_2_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : updatedEntry_2_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : updatedEntry_2_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : updatedEntry_2_uop_aluOp_string = "sra_1";
      ALUOp_passa : updatedEntry_2_uop_aluOp_string = "passa";
      ALUOp_passb : updatedEntry_2_uop_aluOp_string = "passb";
      default : updatedEntry_2_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_uop_bruOp)
      BRUOp_nop : updatedEntry_2_uop_bruOp_string = "nop  ";
      BRUOp_add : updatedEntry_2_uop_bruOp_string = "add  ";
      BRUOp_cadd : updatedEntry_2_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : updatedEntry_2_uop_bruOp_string = "ncadd";
      default : updatedEntry_2_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_roop_aluROOp)
      ALUROOp_reg_1 : updatedEntry_2_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : updatedEntry_2_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : updatedEntry_2_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : updatedEntry_2_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : updatedEntry_2_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : updatedEntry_2_roop_aluROOp_string = "linkreg";
      default : updatedEntry_2_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_roop_cruROOp)
      CRUROOp_id : updatedEntry_2_roop_cruROOp_string = "id";
      CRUROOp_lo : updatedEntry_2_roop_cruROOp_string = "lo";
      CRUROOp_hi : updatedEntry_2_roop_cruROOp_string = "hi";
      default : updatedEntry_2_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_uop_aluOp)
      ALUOp_add : updatedEntry_3_uop_aluOp_string = "add  ";
      ALUOp_sub : updatedEntry_3_uop_aluOp_string = "sub  ";
      ALUOp_slt : updatedEntry_3_uop_aluOp_string = "slt  ";
      ALUOp_sltu : updatedEntry_3_uop_aluOp_string = "sltu ";
      ALUOp_eq : updatedEntry_3_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : updatedEntry_3_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : updatedEntry_3_uop_aluOp_string = "and_1";
      ALUOp_or_1 : updatedEntry_3_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : updatedEntry_3_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : updatedEntry_3_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : updatedEntry_3_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : updatedEntry_3_uop_aluOp_string = "sra_1";
      ALUOp_passa : updatedEntry_3_uop_aluOp_string = "passa";
      ALUOp_passb : updatedEntry_3_uop_aluOp_string = "passb";
      default : updatedEntry_3_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_uop_bruOp)
      BRUOp_nop : updatedEntry_3_uop_bruOp_string = "nop  ";
      BRUOp_add : updatedEntry_3_uop_bruOp_string = "add  ";
      BRUOp_cadd : updatedEntry_3_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : updatedEntry_3_uop_bruOp_string = "ncadd";
      default : updatedEntry_3_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_roop_aluROOp)
      ALUROOp_reg_1 : updatedEntry_3_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : updatedEntry_3_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : updatedEntry_3_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : updatedEntry_3_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : updatedEntry_3_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : updatedEntry_3_roop_aluROOp_string = "linkreg";
      default : updatedEntry_3_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_roop_cruROOp)
      CRUROOp_id : updatedEntry_3_roop_cruROOp_string = "id";
      CRUROOp_lo : updatedEntry_3_roop_cruROOp_string = "lo";
      CRUROOp_hi : updatedEntry_3_roop_cruROOp_string = "hi";
      default : updatedEntry_3_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(appendEntry_uop_aluOp)
      ALUOp_add : appendEntry_uop_aluOp_string = "add  ";
      ALUOp_sub : appendEntry_uop_aluOp_string = "sub  ";
      ALUOp_slt : appendEntry_uop_aluOp_string = "slt  ";
      ALUOp_sltu : appendEntry_uop_aluOp_string = "sltu ";
      ALUOp_eq : appendEntry_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : appendEntry_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : appendEntry_uop_aluOp_string = "and_1";
      ALUOp_or_1 : appendEntry_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : appendEntry_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : appendEntry_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : appendEntry_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : appendEntry_uop_aluOp_string = "sra_1";
      ALUOp_passa : appendEntry_uop_aluOp_string = "passa";
      ALUOp_passb : appendEntry_uop_aluOp_string = "passb";
      default : appendEntry_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(appendEntry_uop_bruOp)
      BRUOp_nop : appendEntry_uop_bruOp_string = "nop  ";
      BRUOp_add : appendEntry_uop_bruOp_string = "add  ";
      BRUOp_cadd : appendEntry_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : appendEntry_uop_bruOp_string = "ncadd";
      default : appendEntry_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(appendEntry_roop_aluROOp)
      ALUROOp_reg_1 : appendEntry_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : appendEntry_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : appendEntry_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : appendEntry_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : appendEntry_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : appendEntry_roop_aluROOp_string = "linkreg";
      default : appendEntry_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(appendEntry_roop_cruROOp)
      CRUROOp_id : appendEntry_roop_cruROOp_string = "id";
      CRUROOp_lo : appendEntry_roop_cruROOp_string = "lo";
      CRUROOp_hi : appendEntry_roop_cruROOp_string = "hi";
      default : appendEntry_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(queueNext_0_uop_aluOp)
      ALUOp_add : queueNext_0_uop_aluOp_string = "add  ";
      ALUOp_sub : queueNext_0_uop_aluOp_string = "sub  ";
      ALUOp_slt : queueNext_0_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queueNext_0_uop_aluOp_string = "sltu ";
      ALUOp_eq : queueNext_0_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queueNext_0_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queueNext_0_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queueNext_0_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queueNext_0_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queueNext_0_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queueNext_0_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queueNext_0_uop_aluOp_string = "sra_1";
      ALUOp_passa : queueNext_0_uop_aluOp_string = "passa";
      ALUOp_passb : queueNext_0_uop_aluOp_string = "passb";
      default : queueNext_0_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_0_uop_bruOp)
      BRUOp_nop : queueNext_0_uop_bruOp_string = "nop  ";
      BRUOp_add : queueNext_0_uop_bruOp_string = "add  ";
      BRUOp_cadd : queueNext_0_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queueNext_0_uop_bruOp_string = "ncadd";
      default : queueNext_0_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_0_roop_aluROOp)
      ALUROOp_reg_1 : queueNext_0_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queueNext_0_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queueNext_0_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queueNext_0_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queueNext_0_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queueNext_0_roop_aluROOp_string = "linkreg";
      default : queueNext_0_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_0_roop_cruROOp)
      CRUROOp_id : queueNext_0_roop_cruROOp_string = "id";
      CRUROOp_lo : queueNext_0_roop_cruROOp_string = "lo";
      CRUROOp_hi : queueNext_0_roop_cruROOp_string = "hi";
      default : queueNext_0_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(queueNext_1_uop_aluOp)
      ALUOp_add : queueNext_1_uop_aluOp_string = "add  ";
      ALUOp_sub : queueNext_1_uop_aluOp_string = "sub  ";
      ALUOp_slt : queueNext_1_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queueNext_1_uop_aluOp_string = "sltu ";
      ALUOp_eq : queueNext_1_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queueNext_1_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queueNext_1_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queueNext_1_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queueNext_1_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queueNext_1_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queueNext_1_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queueNext_1_uop_aluOp_string = "sra_1";
      ALUOp_passa : queueNext_1_uop_aluOp_string = "passa";
      ALUOp_passb : queueNext_1_uop_aluOp_string = "passb";
      default : queueNext_1_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_1_uop_bruOp)
      BRUOp_nop : queueNext_1_uop_bruOp_string = "nop  ";
      BRUOp_add : queueNext_1_uop_bruOp_string = "add  ";
      BRUOp_cadd : queueNext_1_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queueNext_1_uop_bruOp_string = "ncadd";
      default : queueNext_1_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_1_roop_aluROOp)
      ALUROOp_reg_1 : queueNext_1_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queueNext_1_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queueNext_1_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queueNext_1_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queueNext_1_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queueNext_1_roop_aluROOp_string = "linkreg";
      default : queueNext_1_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_1_roop_cruROOp)
      CRUROOp_id : queueNext_1_roop_cruROOp_string = "id";
      CRUROOp_lo : queueNext_1_roop_cruROOp_string = "lo";
      CRUROOp_hi : queueNext_1_roop_cruROOp_string = "hi";
      default : queueNext_1_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(queueNext_2_uop_aluOp)
      ALUOp_add : queueNext_2_uop_aluOp_string = "add  ";
      ALUOp_sub : queueNext_2_uop_aluOp_string = "sub  ";
      ALUOp_slt : queueNext_2_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queueNext_2_uop_aluOp_string = "sltu ";
      ALUOp_eq : queueNext_2_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queueNext_2_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queueNext_2_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queueNext_2_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queueNext_2_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queueNext_2_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queueNext_2_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queueNext_2_uop_aluOp_string = "sra_1";
      ALUOp_passa : queueNext_2_uop_aluOp_string = "passa";
      ALUOp_passb : queueNext_2_uop_aluOp_string = "passb";
      default : queueNext_2_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_2_uop_bruOp)
      BRUOp_nop : queueNext_2_uop_bruOp_string = "nop  ";
      BRUOp_add : queueNext_2_uop_bruOp_string = "add  ";
      BRUOp_cadd : queueNext_2_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queueNext_2_uop_bruOp_string = "ncadd";
      default : queueNext_2_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_2_roop_aluROOp)
      ALUROOp_reg_1 : queueNext_2_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queueNext_2_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queueNext_2_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queueNext_2_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queueNext_2_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queueNext_2_roop_aluROOp_string = "linkreg";
      default : queueNext_2_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_2_roop_cruROOp)
      CRUROOp_id : queueNext_2_roop_cruROOp_string = "id";
      CRUROOp_lo : queueNext_2_roop_cruROOp_string = "lo";
      CRUROOp_hi : queueNext_2_roop_cruROOp_string = "hi";
      default : queueNext_2_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(queueNext_3_uop_aluOp)
      ALUOp_add : queueNext_3_uop_aluOp_string = "add  ";
      ALUOp_sub : queueNext_3_uop_aluOp_string = "sub  ";
      ALUOp_slt : queueNext_3_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queueNext_3_uop_aluOp_string = "sltu ";
      ALUOp_eq : queueNext_3_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queueNext_3_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queueNext_3_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queueNext_3_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queueNext_3_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queueNext_3_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queueNext_3_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queueNext_3_uop_aluOp_string = "sra_1";
      ALUOp_passa : queueNext_3_uop_aluOp_string = "passa";
      ALUOp_passb : queueNext_3_uop_aluOp_string = "passb";
      default : queueNext_3_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_3_uop_bruOp)
      BRUOp_nop : queueNext_3_uop_bruOp_string = "nop  ";
      BRUOp_add : queueNext_3_uop_bruOp_string = "add  ";
      BRUOp_cadd : queueNext_3_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queueNext_3_uop_bruOp_string = "ncadd";
      default : queueNext_3_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_3_roop_aluROOp)
      ALUROOp_reg_1 : queueNext_3_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queueNext_3_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queueNext_3_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queueNext_3_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queueNext_3_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queueNext_3_roop_aluROOp_string = "linkreg";
      default : queueNext_3_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_3_roop_cruROOp)
      CRUROOp_id : queueNext_3_roop_cruROOp_string = "id";
      CRUROOp_lo : queueNext_3_roop_cruROOp_string = "lo";
      CRUROOp_hi : queueNext_3_roop_cruROOp_string = "hi";
      default : queueNext_3_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(issueEntry_uop_aluOp)
      ALUOp_add : issueEntry_uop_aluOp_string = "add  ";
      ALUOp_sub : issueEntry_uop_aluOp_string = "sub  ";
      ALUOp_slt : issueEntry_uop_aluOp_string = "slt  ";
      ALUOp_sltu : issueEntry_uop_aluOp_string = "sltu ";
      ALUOp_eq : issueEntry_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : issueEntry_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : issueEntry_uop_aluOp_string = "and_1";
      ALUOp_or_1 : issueEntry_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : issueEntry_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : issueEntry_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : issueEntry_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : issueEntry_uop_aluOp_string = "sra_1";
      ALUOp_passa : issueEntry_uop_aluOp_string = "passa";
      ALUOp_passb : issueEntry_uop_aluOp_string = "passb";
      default : issueEntry_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(issueEntry_uop_bruOp)
      BRUOp_nop : issueEntry_uop_bruOp_string = "nop  ";
      BRUOp_add : issueEntry_uop_bruOp_string = "add  ";
      BRUOp_cadd : issueEntry_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : issueEntry_uop_bruOp_string = "ncadd";
      default : issueEntry_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(issueEntry_roop_aluROOp)
      ALUROOp_reg_1 : issueEntry_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : issueEntry_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : issueEntry_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : issueEntry_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : issueEntry_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : issueEntry_roop_aluROOp_string = "linkreg";
      default : issueEntry_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(issueEntry_roop_cruROOp)
      CRUROOp_id : issueEntry_roop_cruROOp_string = "id";
      CRUROOp_lo : issueEntry_roop_cruROOp_string = "lo";
      CRUROOp_hi : issueEntry_roop_cruROOp_string = "hi";
      default : issueEntry_roop_cruROOp_string = "??";
    endcase
  end
  `endif

  always @(*) begin
    readyToIssue[0] = ((queue_0_valid && queue_0_srcReady_0) && queue_0_srcReady_1);
    readyToIssue[1] = ((queue_1_valid && queue_1_srcReady_0) && queue_1_srcReady_1);
    readyToIssue[2] = ((queue_2_valid && queue_2_srcReady_0) && queue_2_srcReady_1);
    readyToIssue[3] = ((queue_3_valid && queue_3_srcReady_0) && queue_3_srcReady_1);
  end

  assign readyToIssue_ohFirst_input = readyToIssue;
  assign readyToIssue_ohFirst_masked = (readyToIssue_ohFirst_input & (~ _zz_readyToIssue_ohFirst_masked));
  assign issueVector = readyToIssue_ohFirst_masked;
  always @(*) begin
    emptyEntry[0] = (! queue_0_valid);
    emptyEntry[1] = (! queue_1_valid);
    emptyEntry[2] = (! queue_2_valid);
    emptyEntry[3] = (! queue_3_valid);
    emptyEntry[4] = 1'b1;
    emptyEntry[0] = (! queue_0_valid);
    emptyEntry[1] = (! queue_1_valid);
    emptyEntry[2] = (! queue_2_valid);
    emptyEntry[3] = (! queue_3_valid);
  end

  assign emptyEntry_ohFirst_input = emptyEntry;
  assign emptyEntry_ohFirst_masked = (emptyEntry_ohFirst_input & (~ _zz_emptyEntry_ohFirst_masked));
  assign writeVector = emptyEntry_ohFirst_masked;
  assign appendEntry_valid = io_input_valid;
  assign appendEntry_robIdx = io_input_payload_robIdx;
  assign appendEntry_branchInfo_predictPC = io_input_payload_branchInfo_predictPC;
  assign appendEntry_branchInfo_predictResult = io_input_payload_branchInfo_predictResult;
  assign appendEntry_exceptionInfo_exception = io_input_payload_exceptionInfo_exception;
  assign appendEntry_exceptionInfo_eCode = io_input_payload_exceptionInfo_eCode;
  assign appendEntry_exceptionInfo_eSubCode = io_input_payload_exceptionInfo_eSubCode;
  assign appendEntry_pc = io_input_payload_pc;
  assign appendEntry_prd = io_input_payload_prd;
  assign appendEntry_psrc_0 = io_input_payload_psrc_0;
  assign appendEntry_psrc_1 = io_input_payload_psrc_1;
  assign appendEntry_imm = io_input_payload_imm;
  assign appendEntry_uop_aluOp = io_input_payload_uop_aluOp;
  assign appendEntry_uop_bruOp = io_input_payload_uop_bruOp;
  assign appendEntry_roop_aluROOp = io_input_payload_roop_aluROOp;
  assign appendEntry_roop_cruROOp = io_input_payload_roop_cruROOp;
  assign appendEntry_srcReady_0 = ((io_input_payload_srcReady_0 || (|{(io_input_payload_psrc_0 == io_writebackSignal_4),{_zz_appendEntry_srcReady_0,{_zz_appendEntry_srcReady_0_1,_zz_appendEntry_srcReady_0_2}}})) || ((|{(_zz_appendEntry_srcReady_0_3 && io_earlyWakeup_7_valid),{_zz_appendEntry_srcReady_0_4,{_zz_appendEntry_srcReady_0_5,_zz_appendEntry_srcReady_0_6}}}) || ((io_input_payload_psrc_0 == io_wakeOut_payload) && io_wakeOut_valid)));
  assign appendEntry_srcReady_1 = ((io_input_payload_srcReady_1 || (|{(io_input_payload_psrc_1 == io_writebackSignal_4),{(io_input_payload_psrc_1 == io_writebackSignal_3),{_zz_appendEntry_srcReady_1,{_zz_appendEntry_srcReady_1_1,_zz_appendEntry_srcReady_1_2}}}})) || ((|{((io_input_payload_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_appendEntry_srcReady_1_3 && io_earlyWakeup_6_valid),{_zz_appendEntry_srcReady_1_4,{_zz_appendEntry_srcReady_1_5,_zz_appendEntry_srcReady_1_6}}}}) || ((io_input_payload_psrc_1 == io_wakeOut_payload) && io_wakeOut_valid)));
  assign updatedEntry_0_valid = queue_0_valid;
  assign updatedEntry_0_robIdx = queue_0_robIdx;
  assign updatedEntry_0_branchInfo_predictPC = queue_0_branchInfo_predictPC;
  assign updatedEntry_0_branchInfo_predictResult = queue_0_branchInfo_predictResult;
  assign updatedEntry_0_exceptionInfo_exception = queue_0_exceptionInfo_exception;
  assign updatedEntry_0_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
  assign updatedEntry_0_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
  assign updatedEntry_0_pc = queue_0_pc;
  assign updatedEntry_0_prd = queue_0_prd;
  assign updatedEntry_0_psrc_0 = queue_0_psrc_0;
  assign updatedEntry_0_psrc_1 = queue_0_psrc_1;
  assign updatedEntry_0_imm = queue_0_imm;
  assign updatedEntry_0_uop_aluOp = queue_0_uop_aluOp;
  assign updatedEntry_0_uop_bruOp = queue_0_uop_bruOp;
  assign updatedEntry_0_roop_aluROOp = queue_0_roop_aluROOp;
  assign updatedEntry_0_roop_cruROOp = queue_0_roop_cruROOp;
  always @(*) begin
    updatedEntry_0_srcReady_0 = queue_0_srcReady_0;
    updatedEntry_0_srcReady_0 = ((queue_0_srcReady_0 || (|{(queue_0_psrc_0 == io_writebackSignal_4),{(queue_0_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_0_srcReady_0,{_zz_updatedEntry_0_srcReady_0_1,_zz_updatedEntry_0_srcReady_0_2}}}})) || ((|{((queue_0_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_0_srcReady_0_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_0_srcReady_0_4,{_zz_updatedEntry_0_srcReady_0_5,_zz_updatedEntry_0_srcReady_0_6}}}}) || ((queue_0_psrc_0 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  always @(*) begin
    updatedEntry_0_srcReady_1 = queue_0_srcReady_1;
    updatedEntry_0_srcReady_1 = ((queue_0_srcReady_1 || (|{(queue_0_psrc_1 == io_writebackSignal_4),{(queue_0_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_0_srcReady_1,{_zz_updatedEntry_0_srcReady_1_1,_zz_updatedEntry_0_srcReady_1_2}}}})) || ((|{((queue_0_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_0_srcReady_1_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_0_srcReady_1_4,{_zz_updatedEntry_0_srcReady_1_5,_zz_updatedEntry_0_srcReady_1_6}}}}) || ((queue_0_psrc_1 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  assign updatedEntry_1_valid = queue_1_valid;
  assign updatedEntry_1_robIdx = queue_1_robIdx;
  assign updatedEntry_1_branchInfo_predictPC = queue_1_branchInfo_predictPC;
  assign updatedEntry_1_branchInfo_predictResult = queue_1_branchInfo_predictResult;
  assign updatedEntry_1_exceptionInfo_exception = queue_1_exceptionInfo_exception;
  assign updatedEntry_1_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
  assign updatedEntry_1_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
  assign updatedEntry_1_pc = queue_1_pc;
  assign updatedEntry_1_prd = queue_1_prd;
  assign updatedEntry_1_psrc_0 = queue_1_psrc_0;
  assign updatedEntry_1_psrc_1 = queue_1_psrc_1;
  assign updatedEntry_1_imm = queue_1_imm;
  assign updatedEntry_1_uop_aluOp = queue_1_uop_aluOp;
  assign updatedEntry_1_uop_bruOp = queue_1_uop_bruOp;
  assign updatedEntry_1_roop_aluROOp = queue_1_roop_aluROOp;
  assign updatedEntry_1_roop_cruROOp = queue_1_roop_cruROOp;
  always @(*) begin
    updatedEntry_1_srcReady_0 = queue_1_srcReady_0;
    updatedEntry_1_srcReady_0 = ((queue_1_srcReady_0 || (|{(queue_1_psrc_0 == io_writebackSignal_4),{(queue_1_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_1_srcReady_0,{_zz_updatedEntry_1_srcReady_0_1,_zz_updatedEntry_1_srcReady_0_2}}}})) || ((|{((queue_1_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_1_srcReady_0_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_1_srcReady_0_4,{_zz_updatedEntry_1_srcReady_0_5,_zz_updatedEntry_1_srcReady_0_6}}}}) || ((queue_1_psrc_0 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  always @(*) begin
    updatedEntry_1_srcReady_1 = queue_1_srcReady_1;
    updatedEntry_1_srcReady_1 = ((queue_1_srcReady_1 || (|{(queue_1_psrc_1 == io_writebackSignal_4),{(queue_1_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_1_srcReady_1,{_zz_updatedEntry_1_srcReady_1_1,_zz_updatedEntry_1_srcReady_1_2}}}})) || ((|{((queue_1_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_1_srcReady_1_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_1_srcReady_1_4,{_zz_updatedEntry_1_srcReady_1_5,_zz_updatedEntry_1_srcReady_1_6}}}}) || ((queue_1_psrc_1 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  assign updatedEntry_2_valid = queue_2_valid;
  assign updatedEntry_2_robIdx = queue_2_robIdx;
  assign updatedEntry_2_branchInfo_predictPC = queue_2_branchInfo_predictPC;
  assign updatedEntry_2_branchInfo_predictResult = queue_2_branchInfo_predictResult;
  assign updatedEntry_2_exceptionInfo_exception = queue_2_exceptionInfo_exception;
  assign updatedEntry_2_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
  assign updatedEntry_2_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
  assign updatedEntry_2_pc = queue_2_pc;
  assign updatedEntry_2_prd = queue_2_prd;
  assign updatedEntry_2_psrc_0 = queue_2_psrc_0;
  assign updatedEntry_2_psrc_1 = queue_2_psrc_1;
  assign updatedEntry_2_imm = queue_2_imm;
  assign updatedEntry_2_uop_aluOp = queue_2_uop_aluOp;
  assign updatedEntry_2_uop_bruOp = queue_2_uop_bruOp;
  assign updatedEntry_2_roop_aluROOp = queue_2_roop_aluROOp;
  assign updatedEntry_2_roop_cruROOp = queue_2_roop_cruROOp;
  always @(*) begin
    updatedEntry_2_srcReady_0 = queue_2_srcReady_0;
    updatedEntry_2_srcReady_0 = ((queue_2_srcReady_0 || (|{(queue_2_psrc_0 == io_writebackSignal_4),{(queue_2_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_2_srcReady_0,{_zz_updatedEntry_2_srcReady_0_1,_zz_updatedEntry_2_srcReady_0_2}}}})) || ((|{((queue_2_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_2_srcReady_0_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_2_srcReady_0_4,{_zz_updatedEntry_2_srcReady_0_5,_zz_updatedEntry_2_srcReady_0_6}}}}) || ((queue_2_psrc_0 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  always @(*) begin
    updatedEntry_2_srcReady_1 = queue_2_srcReady_1;
    updatedEntry_2_srcReady_1 = ((queue_2_srcReady_1 || (|{(queue_2_psrc_1 == io_writebackSignal_4),{(queue_2_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_2_srcReady_1,{_zz_updatedEntry_2_srcReady_1_1,_zz_updatedEntry_2_srcReady_1_2}}}})) || ((|{((queue_2_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_2_srcReady_1_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_2_srcReady_1_4,{_zz_updatedEntry_2_srcReady_1_5,_zz_updatedEntry_2_srcReady_1_6}}}}) || ((queue_2_psrc_1 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  assign updatedEntry_3_valid = queue_3_valid;
  assign updatedEntry_3_robIdx = queue_3_robIdx;
  assign updatedEntry_3_branchInfo_predictPC = queue_3_branchInfo_predictPC;
  assign updatedEntry_3_branchInfo_predictResult = queue_3_branchInfo_predictResult;
  assign updatedEntry_3_exceptionInfo_exception = queue_3_exceptionInfo_exception;
  assign updatedEntry_3_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
  assign updatedEntry_3_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
  assign updatedEntry_3_pc = queue_3_pc;
  assign updatedEntry_3_prd = queue_3_prd;
  assign updatedEntry_3_psrc_0 = queue_3_psrc_0;
  assign updatedEntry_3_psrc_1 = queue_3_psrc_1;
  assign updatedEntry_3_imm = queue_3_imm;
  assign updatedEntry_3_uop_aluOp = queue_3_uop_aluOp;
  assign updatedEntry_3_uop_bruOp = queue_3_uop_bruOp;
  assign updatedEntry_3_roop_aluROOp = queue_3_roop_aluROOp;
  assign updatedEntry_3_roop_cruROOp = queue_3_roop_cruROOp;
  always @(*) begin
    updatedEntry_3_srcReady_0 = queue_3_srcReady_0;
    updatedEntry_3_srcReady_0 = ((queue_3_srcReady_0 || (|{(queue_3_psrc_0 == io_writebackSignal_4),{(queue_3_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_3_srcReady_0,{_zz_updatedEntry_3_srcReady_0_1,_zz_updatedEntry_3_srcReady_0_2}}}})) || ((|{((queue_3_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_3_srcReady_0_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_3_srcReady_0_4,{_zz_updatedEntry_3_srcReady_0_5,_zz_updatedEntry_3_srcReady_0_6}}}}) || ((queue_3_psrc_0 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  always @(*) begin
    updatedEntry_3_srcReady_1 = queue_3_srcReady_1;
    updatedEntry_3_srcReady_1 = ((queue_3_srcReady_1 || (|{(queue_3_psrc_1 == io_writebackSignal_4),{(queue_3_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_3_srcReady_1,{_zz_updatedEntry_3_srcReady_1_1,_zz_updatedEntry_3_srcReady_1_2}}}})) || ((|{((queue_3_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_3_srcReady_1_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_3_srcReady_1_4,{_zz_updatedEntry_3_srcReady_1_5,_zz_updatedEntry_3_srcReady_1_6}}}}) || ((queue_3_psrc_1 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  always @(*) begin
    shiftAhead[0] = ((|readyToIssue[0 : 0]) && io_output_ready);
    shiftAhead[1] = ((|readyToIssue[1 : 0]) && io_output_ready);
    shiftAhead[2] = ((|readyToIssue[2 : 0]) && io_output_ready);
    shiftAhead[3] = ((|readyToIssue[3 : 0]) && io_output_ready);
  end

  assign when_IssueQueue_l81 = shiftAhead[0];
  assign when_IssueQueue_l83 = writeVector[1];
  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_valid = appendEntry_valid;
      end else begin
        queueNext_0_valid = queue_1_valid;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_valid = appendEntry_valid;
      end else begin
        queueNext_0_valid = queue_0_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_0_robIdx = queue_1_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_0_robIdx = queue_0_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_0_branchInfo_predictPC = queue_1_branchInfo_predictPC;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_0_branchInfo_predictPC = queue_0_branchInfo_predictPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_0_branchInfo_predictResult = queue_1_branchInfo_predictResult;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_0_branchInfo_predictResult = queue_0_branchInfo_predictResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_0_exceptionInfo_exception = queue_1_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_0_exceptionInfo_exception = queue_0_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_0_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_0_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_0_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_0_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_pc = appendEntry_pc;
      end else begin
        queueNext_0_pc = queue_1_pc;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_pc = appendEntry_pc;
      end else begin
        queueNext_0_pc = queue_0_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_prd = appendEntry_prd;
      end else begin
        queueNext_0_prd = queue_1_prd;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_prd = appendEntry_prd;
      end else begin
        queueNext_0_prd = queue_0_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_0_psrc_0 = queue_1_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_0_psrc_0 = queue_0_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_0_psrc_1 = queue_1_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_0_psrc_1 = queue_0_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_imm = appendEntry_imm;
      end else begin
        queueNext_0_imm = queue_1_imm;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_imm = appendEntry_imm;
      end else begin
        queueNext_0_imm = queue_0_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_0_uop_aluOp = queue_1_uop_aluOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_0_uop_aluOp = queue_0_uop_aluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_0_uop_bruOp = queue_1_uop_bruOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_0_uop_bruOp = queue_0_uop_bruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_0_roop_aluROOp = queue_1_roop_aluROOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_0_roop_aluROOp = queue_0_roop_aluROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_roop_cruROOp = appendEntry_roop_cruROOp;
      end else begin
        queueNext_0_roop_cruROOp = queue_1_roop_cruROOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_roop_cruROOp = appendEntry_roop_cruROOp;
      end else begin
        queueNext_0_roop_cruROOp = queue_0_roop_cruROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_0_srcReady_0 = queue_1_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_0_srcReady_0 = queue_0_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_0_srcReady_1 = queue_1_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_0_srcReady_1 = queue_0_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96 = writeVector[0];
  assign when_IssueQueue_l81_1 = shiftAhead[1];
  assign when_IssueQueue_l83_1 = writeVector[2];
  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_valid = appendEntry_valid;
      end else begin
        queueNext_1_valid = queue_2_valid;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_valid = appendEntry_valid;
      end else begin
        queueNext_1_valid = queue_1_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_1_robIdx = queue_2_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_1_robIdx = queue_1_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_1_branchInfo_predictPC = queue_2_branchInfo_predictPC;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_1_branchInfo_predictPC = queue_1_branchInfo_predictPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_1_branchInfo_predictResult = queue_2_branchInfo_predictResult;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_1_branchInfo_predictResult = queue_1_branchInfo_predictResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_1_exceptionInfo_exception = queue_2_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_1_exceptionInfo_exception = queue_1_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_1_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_1_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_1_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_1_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_pc = appendEntry_pc;
      end else begin
        queueNext_1_pc = queue_2_pc;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_pc = appendEntry_pc;
      end else begin
        queueNext_1_pc = queue_1_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_prd = appendEntry_prd;
      end else begin
        queueNext_1_prd = queue_2_prd;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_prd = appendEntry_prd;
      end else begin
        queueNext_1_prd = queue_1_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_1_psrc_0 = queue_2_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_1_psrc_0 = queue_1_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_1_psrc_1 = queue_2_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_1_psrc_1 = queue_1_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_imm = appendEntry_imm;
      end else begin
        queueNext_1_imm = queue_2_imm;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_imm = appendEntry_imm;
      end else begin
        queueNext_1_imm = queue_1_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_1_uop_aluOp = queue_2_uop_aluOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_1_uop_aluOp = queue_1_uop_aluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_1_uop_bruOp = queue_2_uop_bruOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_1_uop_bruOp = queue_1_uop_bruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_1_roop_aluROOp = queue_2_roop_aluROOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_1_roop_aluROOp = queue_1_roop_aluROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_roop_cruROOp = appendEntry_roop_cruROOp;
      end else begin
        queueNext_1_roop_cruROOp = queue_2_roop_cruROOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_roop_cruROOp = appendEntry_roop_cruROOp;
      end else begin
        queueNext_1_roop_cruROOp = queue_1_roop_cruROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_1_srcReady_0 = queue_2_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_1_srcReady_0 = queue_1_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_1_srcReady_1 = queue_2_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_1_srcReady_1 = queue_1_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_1 = writeVector[1];
  assign when_IssueQueue_l81_2 = shiftAhead[2];
  assign when_IssueQueue_l83_2 = writeVector[3];
  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_valid = appendEntry_valid;
      end else begin
        queueNext_2_valid = queue_3_valid;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_valid = appendEntry_valid;
      end else begin
        queueNext_2_valid = queue_2_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_2_robIdx = queue_3_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_2_robIdx = queue_2_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_2_branchInfo_predictPC = queue_3_branchInfo_predictPC;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_2_branchInfo_predictPC = queue_2_branchInfo_predictPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_2_branchInfo_predictResult = queue_3_branchInfo_predictResult;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_2_branchInfo_predictResult = queue_2_branchInfo_predictResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_2_exceptionInfo_exception = queue_3_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_2_exceptionInfo_exception = queue_2_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_2_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_2_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_2_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_2_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_pc = appendEntry_pc;
      end else begin
        queueNext_2_pc = queue_3_pc;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_pc = appendEntry_pc;
      end else begin
        queueNext_2_pc = queue_2_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_prd = appendEntry_prd;
      end else begin
        queueNext_2_prd = queue_3_prd;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_prd = appendEntry_prd;
      end else begin
        queueNext_2_prd = queue_2_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_2_psrc_0 = queue_3_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_2_psrc_0 = queue_2_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_2_psrc_1 = queue_3_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_2_psrc_1 = queue_2_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_imm = appendEntry_imm;
      end else begin
        queueNext_2_imm = queue_3_imm;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_imm = appendEntry_imm;
      end else begin
        queueNext_2_imm = queue_2_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_2_uop_aluOp = queue_3_uop_aluOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_2_uop_aluOp = queue_2_uop_aluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_2_uop_bruOp = queue_3_uop_bruOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_2_uop_bruOp = queue_2_uop_bruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_2_roop_aluROOp = queue_3_roop_aluROOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_2_roop_aluROOp = queue_2_roop_aluROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_roop_cruROOp = appendEntry_roop_cruROOp;
      end else begin
        queueNext_2_roop_cruROOp = queue_3_roop_cruROOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_roop_cruROOp = appendEntry_roop_cruROOp;
      end else begin
        queueNext_2_roop_cruROOp = queue_2_roop_cruROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_2_srcReady_0 = queue_3_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_2_srcReady_0 = queue_2_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_2_srcReady_1 = queue_3_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_2_srcReady_1 = queue_2_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_2 = writeVector[2];
  assign when_IssueQueue_l81_3 = shiftAhead[3];
  assign when_IssueQueue_l89 = writeVector[4];
  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_valid = appendEntry_valid;
      end else begin
        queueNext_3_valid = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_valid = appendEntry_valid;
      end else begin
        queueNext_3_valid = queue_3_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_3_robIdx = 5'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_3_robIdx = queue_3_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_3_branchInfo_predictPC = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_3_branchInfo_predictPC = queue_3_branchInfo_predictPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_3_branchInfo_predictResult = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_3_branchInfo_predictResult = queue_3_branchInfo_predictResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_3_exceptionInfo_exception = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_3_exceptionInfo_exception = queue_3_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_3_exceptionInfo_eCode = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_3_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_3_exceptionInfo_eSubCode = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_3_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_pc = appendEntry_pc;
      end else begin
        queueNext_3_pc = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_pc = appendEntry_pc;
      end else begin
        queueNext_3_pc = queue_3_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_prd = appendEntry_prd;
      end else begin
        queueNext_3_prd = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_prd = appendEntry_prd;
      end else begin
        queueNext_3_prd = queue_3_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_3_psrc_0 = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_3_psrc_0 = queue_3_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_3_psrc_1 = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_3_psrc_1 = queue_3_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_imm = appendEntry_imm;
      end else begin
        queueNext_3_imm = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_imm = appendEntry_imm;
      end else begin
        queueNext_3_imm = queue_3_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_3_uop_aluOp = ALUOp_add;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_3_uop_aluOp = queue_3_uop_aluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_3_uop_bruOp = BRUOp_nop;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_3_uop_bruOp = queue_3_uop_bruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_3_roop_aluROOp = ALUROOp_reg_1;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_3_roop_aluROOp = queue_3_roop_aluROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_roop_cruROOp = appendEntry_roop_cruROOp;
      end else begin
        queueNext_3_roop_cruROOp = CRUROOp_id;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_roop_cruROOp = appendEntry_roop_cruROOp;
      end else begin
        queueNext_3_roop_cruROOp = queue_3_roop_cruROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_3_srcReady_0 = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_3_srcReady_0 = queue_3_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_3_srcReady_1 = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_3_srcReady_1 = queue_3_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_3 = writeVector[3];
  always @(*) begin
    _zz_io_csrInQueue[0] = ((queue_0_roop_aluROOp == ALUROOp_csr) && queue_0_valid);
    _zz_io_csrInQueue[1] = ((queue_1_roop_aluROOp == ALUROOp_csr) && queue_1_valid);
    _zz_io_csrInQueue[2] = ((queue_2_roop_aluROOp == ALUROOp_csr) && queue_2_valid);
    _zz_io_csrInQueue[3] = ((queue_3_roop_aluROOp == ALUROOp_csr) && queue_3_valid);
  end

  assign io_csrInQueue = (|_zz_io_csrInQueue);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_input_ready = ((|emptyEntry[3 : 0]) || io_output_fire);
  assign _zz_issueEntry_valid = issueVector[3];
  assign _zz_issueEntry_valid_1 = (issueVector[1] || _zz_issueEntry_valid);
  assign _zz_issueEntry_valid_2 = (issueVector[2] || _zz_issueEntry_valid);
  assign _zz_issueEntry_valid_3 = {_zz_issueEntry_valid_2,_zz_issueEntry_valid_1};
  assign issueEntry_valid = _zz_issueEntry_valid_4;
  assign issueEntry_robIdx = _zz_issueEntry_robIdx;
  assign issueEntry_branchInfo_predictPC = _zz_issueEntry_branchInfo_predictPC;
  assign issueEntry_branchInfo_predictResult = _zz_issueEntry_branchInfo_predictResult;
  assign issueEntry_exceptionInfo_exception = _zz_issueEntry_exceptionInfo_exception;
  assign issueEntry_exceptionInfo_eCode = _zz_issueEntry_exceptionInfo_eCode;
  assign issueEntry_exceptionInfo_eSubCode = _zz_issueEntry_exceptionInfo_eSubCode;
  assign issueEntry_pc = _zz_issueEntry_pc;
  assign issueEntry_prd = _zz_issueEntry_prd;
  assign issueEntry_psrc_0 = _zz_issueEntry_psrc_0;
  assign issueEntry_psrc_1 = _zz_issueEntry_psrc_1;
  assign issueEntry_imm = _zz_issueEntry_imm;
  assign issueEntry_uop_aluOp = _zz_issueEntry_uop_aluOp;
  assign issueEntry_uop_bruOp = _zz_issueEntry_uop_bruOp;
  assign issueEntry_roop_aluROOp = _zz_issueEntry_roop_aluROOp;
  assign issueEntry_roop_cruROOp = _zz_issueEntry_roop_cruROOp;
  assign issueEntry_srcReady_0 = _zz_issueEntry_srcReady_0;
  assign issueEntry_srcReady_1 = _zz_issueEntry_srcReady_1;
  assign io_output_valid = (|readyToIssue);
  assign io_output_payload_robIdx = issueEntry_robIdx;
  assign io_output_payload_branchInfo_predictPC = issueEntry_branchInfo_predictPC;
  assign io_output_payload_branchInfo_predictResult = issueEntry_branchInfo_predictResult;
  assign io_output_payload_exceptionInfo_exception = issueEntry_exceptionInfo_exception;
  assign io_output_payload_exceptionInfo_eCode = issueEntry_exceptionInfo_eCode;
  assign io_output_payload_exceptionInfo_eSubCode = issueEntry_exceptionInfo_eSubCode;
  assign io_output_payload_pc = issueEntry_pc;
  assign io_output_payload_prd = issueEntry_prd;
  assign io_output_payload_psrc_0 = issueEntry_psrc_0;
  assign io_output_payload_psrc_1 = issueEntry_psrc_1;
  assign io_output_payload_imm = issueEntry_imm;
  assign io_output_payload_uop_aluOp = issueEntry_uop_aluOp;
  assign io_output_payload_uop_bruOp = issueEntry_uop_bruOp;
  assign io_output_payload_roop_aluROOp = issueEntry_roop_aluROOp;
  assign io_output_payload_roop_cruROOp = issueEntry_roop_cruROOp;
  assign io_wakeOut_payload = issueEntry_prd;
  assign io_wakeOut_valid = io_output_fire;
  always @(posedge aclk) begin
    if(!cpuClockingArea_areaFlushReset_newReset) begin
      queue_0_valid <= 1'b0;
      queue_0_robIdx <= 5'h00;
      queue_0_branchInfo_predictPC <= 32'h00000000;
      queue_0_branchInfo_predictResult <= 1'b0;
      queue_0_exceptionInfo_exception <= 1'b0;
      queue_0_exceptionInfo_eCode <= 6'h00;
      queue_0_exceptionInfo_eSubCode <= 1'b0;
      queue_0_pc <= 32'h00000000;
      queue_0_prd <= 6'h00;
      queue_0_psrc_0 <= 6'h00;
      queue_0_psrc_1 <= 6'h00;
      queue_0_imm <= 32'h00000000;
      queue_0_uop_aluOp <= ALUOp_add;
      queue_0_uop_bruOp <= BRUOp_nop;
      queue_0_roop_aluROOp <= ALUROOp_reg_1;
      queue_0_roop_cruROOp <= CRUROOp_id;
      queue_0_srcReady_0 <= 1'b0;
      queue_0_srcReady_1 <= 1'b0;
      queue_1_valid <= 1'b0;
      queue_1_robIdx <= 5'h00;
      queue_1_branchInfo_predictPC <= 32'h00000000;
      queue_1_branchInfo_predictResult <= 1'b0;
      queue_1_exceptionInfo_exception <= 1'b0;
      queue_1_exceptionInfo_eCode <= 6'h00;
      queue_1_exceptionInfo_eSubCode <= 1'b0;
      queue_1_pc <= 32'h00000000;
      queue_1_prd <= 6'h00;
      queue_1_psrc_0 <= 6'h00;
      queue_1_psrc_1 <= 6'h00;
      queue_1_imm <= 32'h00000000;
      queue_1_uop_aluOp <= ALUOp_add;
      queue_1_uop_bruOp <= BRUOp_nop;
      queue_1_roop_aluROOp <= ALUROOp_reg_1;
      queue_1_roop_cruROOp <= CRUROOp_id;
      queue_1_srcReady_0 <= 1'b0;
      queue_1_srcReady_1 <= 1'b0;
      queue_2_valid <= 1'b0;
      queue_2_robIdx <= 5'h00;
      queue_2_branchInfo_predictPC <= 32'h00000000;
      queue_2_branchInfo_predictResult <= 1'b0;
      queue_2_exceptionInfo_exception <= 1'b0;
      queue_2_exceptionInfo_eCode <= 6'h00;
      queue_2_exceptionInfo_eSubCode <= 1'b0;
      queue_2_pc <= 32'h00000000;
      queue_2_prd <= 6'h00;
      queue_2_psrc_0 <= 6'h00;
      queue_2_psrc_1 <= 6'h00;
      queue_2_imm <= 32'h00000000;
      queue_2_uop_aluOp <= ALUOp_add;
      queue_2_uop_bruOp <= BRUOp_nop;
      queue_2_roop_aluROOp <= ALUROOp_reg_1;
      queue_2_roop_cruROOp <= CRUROOp_id;
      queue_2_srcReady_0 <= 1'b0;
      queue_2_srcReady_1 <= 1'b0;
      queue_3_valid <= 1'b0;
      queue_3_robIdx <= 5'h00;
      queue_3_branchInfo_predictPC <= 32'h00000000;
      queue_3_branchInfo_predictResult <= 1'b0;
      queue_3_exceptionInfo_exception <= 1'b0;
      queue_3_exceptionInfo_eCode <= 6'h00;
      queue_3_exceptionInfo_eSubCode <= 1'b0;
      queue_3_pc <= 32'h00000000;
      queue_3_prd <= 6'h00;
      queue_3_psrc_0 <= 6'h00;
      queue_3_psrc_1 <= 6'h00;
      queue_3_imm <= 32'h00000000;
      queue_3_uop_aluOp <= ALUOp_add;
      queue_3_uop_bruOp <= BRUOp_nop;
      queue_3_roop_aluROOp <= ALUROOp_reg_1;
      queue_3_roop_cruROOp <= CRUROOp_id;
      queue_3_srcReady_0 <= 1'b0;
      queue_3_srcReady_1 <= 1'b0;
    end else begin
      queue_0_valid <= queueNext_0_valid;
      queue_0_robIdx <= queueNext_0_robIdx;
      queue_0_branchInfo_predictPC <= queueNext_0_branchInfo_predictPC;
      queue_0_branchInfo_predictResult <= queueNext_0_branchInfo_predictResult;
      queue_0_exceptionInfo_exception <= queueNext_0_exceptionInfo_exception;
      queue_0_exceptionInfo_eCode <= queueNext_0_exceptionInfo_eCode;
      queue_0_exceptionInfo_eSubCode <= queueNext_0_exceptionInfo_eSubCode;
      queue_0_pc <= queueNext_0_pc;
      queue_0_prd <= queueNext_0_prd;
      queue_0_psrc_0 <= queueNext_0_psrc_0;
      queue_0_psrc_1 <= queueNext_0_psrc_1;
      queue_0_imm <= queueNext_0_imm;
      queue_0_uop_aluOp <= queueNext_0_uop_aluOp;
      queue_0_uop_bruOp <= queueNext_0_uop_bruOp;
      queue_0_roop_aluROOp <= queueNext_0_roop_aluROOp;
      queue_0_roop_cruROOp <= queueNext_0_roop_cruROOp;
      queue_0_srcReady_0 <= queueNext_0_srcReady_0;
      queue_0_srcReady_1 <= queueNext_0_srcReady_1;
      queue_1_valid <= queueNext_1_valid;
      queue_1_robIdx <= queueNext_1_robIdx;
      queue_1_branchInfo_predictPC <= queueNext_1_branchInfo_predictPC;
      queue_1_branchInfo_predictResult <= queueNext_1_branchInfo_predictResult;
      queue_1_exceptionInfo_exception <= queueNext_1_exceptionInfo_exception;
      queue_1_exceptionInfo_eCode <= queueNext_1_exceptionInfo_eCode;
      queue_1_exceptionInfo_eSubCode <= queueNext_1_exceptionInfo_eSubCode;
      queue_1_pc <= queueNext_1_pc;
      queue_1_prd <= queueNext_1_prd;
      queue_1_psrc_0 <= queueNext_1_psrc_0;
      queue_1_psrc_1 <= queueNext_1_psrc_1;
      queue_1_imm <= queueNext_1_imm;
      queue_1_uop_aluOp <= queueNext_1_uop_aluOp;
      queue_1_uop_bruOp <= queueNext_1_uop_bruOp;
      queue_1_roop_aluROOp <= queueNext_1_roop_aluROOp;
      queue_1_roop_cruROOp <= queueNext_1_roop_cruROOp;
      queue_1_srcReady_0 <= queueNext_1_srcReady_0;
      queue_1_srcReady_1 <= queueNext_1_srcReady_1;
      queue_2_valid <= queueNext_2_valid;
      queue_2_robIdx <= queueNext_2_robIdx;
      queue_2_branchInfo_predictPC <= queueNext_2_branchInfo_predictPC;
      queue_2_branchInfo_predictResult <= queueNext_2_branchInfo_predictResult;
      queue_2_exceptionInfo_exception <= queueNext_2_exceptionInfo_exception;
      queue_2_exceptionInfo_eCode <= queueNext_2_exceptionInfo_eCode;
      queue_2_exceptionInfo_eSubCode <= queueNext_2_exceptionInfo_eSubCode;
      queue_2_pc <= queueNext_2_pc;
      queue_2_prd <= queueNext_2_prd;
      queue_2_psrc_0 <= queueNext_2_psrc_0;
      queue_2_psrc_1 <= queueNext_2_psrc_1;
      queue_2_imm <= queueNext_2_imm;
      queue_2_uop_aluOp <= queueNext_2_uop_aluOp;
      queue_2_uop_bruOp <= queueNext_2_uop_bruOp;
      queue_2_roop_aluROOp <= queueNext_2_roop_aluROOp;
      queue_2_roop_cruROOp <= queueNext_2_roop_cruROOp;
      queue_2_srcReady_0 <= queueNext_2_srcReady_0;
      queue_2_srcReady_1 <= queueNext_2_srcReady_1;
      queue_3_valid <= queueNext_3_valid;
      queue_3_robIdx <= queueNext_3_robIdx;
      queue_3_branchInfo_predictPC <= queueNext_3_branchInfo_predictPC;
      queue_3_branchInfo_predictResult <= queueNext_3_branchInfo_predictResult;
      queue_3_exceptionInfo_exception <= queueNext_3_exceptionInfo_exception;
      queue_3_exceptionInfo_eCode <= queueNext_3_exceptionInfo_eCode;
      queue_3_exceptionInfo_eSubCode <= queueNext_3_exceptionInfo_eSubCode;
      queue_3_pc <= queueNext_3_pc;
      queue_3_prd <= queueNext_3_prd;
      queue_3_psrc_0 <= queueNext_3_psrc_0;
      queue_3_psrc_1 <= queueNext_3_psrc_1;
      queue_3_imm <= queueNext_3_imm;
      queue_3_uop_aluOp <= queueNext_3_uop_aluOp;
      queue_3_uop_bruOp <= queueNext_3_uop_bruOp;
      queue_3_roop_aluROOp <= queueNext_3_roop_aluROOp;
      queue_3_roop_cruROOp <= queueNext_3_roop_cruROOp;
      queue_3_srcReady_0 <= queueNext_3_srcReady_0;
      queue_3_srcReady_1 <= queueNext_3_srcReady_1;
    end
  end


endmodule

module IssueQueue (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [4:0]    io_input_payload_robIdx,
  input  wire [31:0]   io_input_payload_branchInfo_predictPC,
  input  wire          io_input_payload_branchInfo_predictResult,
  input  wire          io_input_payload_exceptionInfo_exception,
  input  wire [5:0]    io_input_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_input_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_payload_pc,
  input  wire [5:0]    io_input_payload_prd,
  input  wire [5:0]    io_input_payload_psrc_0,
  input  wire [5:0]    io_input_payload_psrc_1,
  input  wire [31:0]   io_input_payload_imm,
  input  wire [3:0]    io_input_payload_uop_aluOp,
  input  wire [1:0]    io_input_payload_uop_bruOp,
  input  wire [1:0]    io_input_payload_uop_cruOp,
  input  wire [2:0]    io_input_payload_roop_aluROOp,
  input  wire          io_input_payload_srcReady_0,
  input  wire          io_input_payload_srcReady_1,
  output wire          io_csrInQueue,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [4:0]    io_output_payload_robIdx,
  output wire [31:0]   io_output_payload_branchInfo_predictPC,
  output wire          io_output_payload_branchInfo_predictResult,
  output wire          io_output_payload_exceptionInfo_exception,
  output wire [5:0]    io_output_payload_exceptionInfo_eCode,
  output wire [0:0]    io_output_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_output_payload_pc,
  output wire [5:0]    io_output_payload_prd,
  output wire [5:0]    io_output_payload_psrc_0,
  output wire [5:0]    io_output_payload_psrc_1,
  output wire [31:0]   io_output_payload_imm,
  output wire [3:0]    io_output_payload_uop_aluOp,
  output wire [1:0]    io_output_payload_uop_bruOp,
  output wire [1:0]    io_output_payload_uop_cruOp,
  output wire [2:0]    io_output_payload_roop_aluROOp,
  input  wire [5:0]    io_writebackSignal_0,
  input  wire [5:0]    io_writebackSignal_1,
  input  wire [5:0]    io_writebackSignal_2,
  input  wire [5:0]    io_writebackSignal_3,
  input  wire [5:0]    io_writebackSignal_4,
  input  wire          io_earlyWakeup_0_valid,
  input  wire [5:0]    io_earlyWakeup_0_payload,
  input  wire          io_earlyWakeup_1_valid,
  input  wire [5:0]    io_earlyWakeup_1_payload,
  input  wire          io_earlyWakeup_2_valid,
  input  wire [5:0]    io_earlyWakeup_2_payload,
  input  wire          io_earlyWakeup_3_valid,
  input  wire [5:0]    io_earlyWakeup_3_payload,
  input  wire          io_earlyWakeup_4_valid,
  input  wire [5:0]    io_earlyWakeup_4_payload,
  input  wire          io_earlyWakeup_5_valid,
  input  wire [5:0]    io_earlyWakeup_5_payload,
  input  wire          io_earlyWakeup_6_valid,
  input  wire [5:0]    io_earlyWakeup_6_payload,
  input  wire          io_earlyWakeup_7_valid,
  input  wire [5:0]    io_earlyWakeup_7_payload,
  output wire          io_wakeOut_valid,
  output wire [5:0]    io_wakeOut_payload,
  input  wire          aclk,
  input  wire          cpuClockingArea_areaFlushReset_newReset
);
  localparam ALUOp_add = 4'd0;
  localparam ALUOp_sub = 4'd1;
  localparam ALUOp_slt = 4'd2;
  localparam ALUOp_sltu = 4'd3;
  localparam ALUOp_eq = 4'd4;
  localparam ALUOp_nor_1 = 4'd5;
  localparam ALUOp_and_1 = 4'd6;
  localparam ALUOp_or_1 = 4'd7;
  localparam ALUOp_xor_1 = 4'd8;
  localparam ALUOp_sll_1 = 4'd9;
  localparam ALUOp_srl_1 = 4'd10;
  localparam ALUOp_sra_1 = 4'd11;
  localparam ALUOp_passa = 4'd12;
  localparam ALUOp_passb = 4'd13;
  localparam BRUOp_nop = 2'd0;
  localparam BRUOp_add = 2'd1;
  localparam BRUOp_cadd = 2'd2;
  localparam BRUOp_ncadd = 2'd3;
  localparam CRUOp_nop = 2'd0;
  localparam CRUOp_pass = 2'd1;
  localparam CRUOp_mask = 2'd2;
  localparam ALUROOp_reg_1 = 3'd0;
  localparam ALUROOp_regimm = 3'd1;
  localparam ALUROOp_pcimm = 3'd2;
  localparam ALUROOp_csr = 3'd3;
  localparam ALUROOp_linkpc = 3'd4;
  localparam ALUROOp_linkreg = 3'd5;

  wire       [3:0]    _zz_readyToIssue_ohFirst_masked;
  wire       [4:0]    _zz_emptyEntry_ohFirst_masked;
  wire                _zz_appendEntry_srcReady_0;
  wire       [0:0]    _zz_appendEntry_srcReady_0_1;
  wire       [1:0]    _zz_appendEntry_srcReady_0_2;
  wire                _zz_appendEntry_srcReady_0_3;
  wire                _zz_appendEntry_srcReady_0_4;
  wire       [0:0]    _zz_appendEntry_srcReady_0_5;
  wire       [4:0]    _zz_appendEntry_srcReady_0_6;
  wire                _zz_appendEntry_srcReady_0_7;
  wire                _zz_appendEntry_srcReady_0_8;
  wire       [0:0]    _zz_appendEntry_srcReady_0_9;
  wire       [0:0]    _zz_appendEntry_srcReady_0_10;
  wire                _zz_appendEntry_srcReady_1;
  wire       [0:0]    _zz_appendEntry_srcReady_1_1;
  wire       [0:0]    _zz_appendEntry_srcReady_1_2;
  wire                _zz_appendEntry_srcReady_1_3;
  wire                _zz_appendEntry_srcReady_1_4;
  wire       [0:0]    _zz_appendEntry_srcReady_1_5;
  wire       [3:0]    _zz_appendEntry_srcReady_1_6;
  wire                _zz_updatedEntry_0_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_0_2;
  wire                _zz_updatedEntry_0_srcReady_0_3;
  wire                _zz_updatedEntry_0_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_0_5;
  wire       [3:0]    _zz_updatedEntry_0_srcReady_0_6;
  wire                _zz_updatedEntry_0_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_1_2;
  wire                _zz_updatedEntry_0_srcReady_1_3;
  wire                _zz_updatedEntry_0_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_0_srcReady_1_5;
  wire       [3:0]    _zz_updatedEntry_0_srcReady_1_6;
  wire                _zz_updatedEntry_1_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_0_2;
  wire                _zz_updatedEntry_1_srcReady_0_3;
  wire                _zz_updatedEntry_1_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_0_5;
  wire       [3:0]    _zz_updatedEntry_1_srcReady_0_6;
  wire                _zz_updatedEntry_1_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_1_2;
  wire                _zz_updatedEntry_1_srcReady_1_3;
  wire                _zz_updatedEntry_1_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_1_srcReady_1_5;
  wire       [3:0]    _zz_updatedEntry_1_srcReady_1_6;
  wire                _zz_updatedEntry_2_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_0_2;
  wire                _zz_updatedEntry_2_srcReady_0_3;
  wire                _zz_updatedEntry_2_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_0_5;
  wire       [3:0]    _zz_updatedEntry_2_srcReady_0_6;
  wire                _zz_updatedEntry_2_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_1_2;
  wire                _zz_updatedEntry_2_srcReady_1_3;
  wire                _zz_updatedEntry_2_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_2_srcReady_1_5;
  wire       [3:0]    _zz_updatedEntry_2_srcReady_1_6;
  wire                _zz_updatedEntry_3_srcReady_0;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_0_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_0_2;
  wire                _zz_updatedEntry_3_srcReady_0_3;
  wire                _zz_updatedEntry_3_srcReady_0_4;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_0_5;
  wire       [3:0]    _zz_updatedEntry_3_srcReady_0_6;
  wire                _zz_updatedEntry_3_srcReady_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_1_1;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_1_2;
  wire                _zz_updatedEntry_3_srcReady_1_3;
  wire                _zz_updatedEntry_3_srcReady_1_4;
  wire       [0:0]    _zz_updatedEntry_3_srcReady_1_5;
  wire       [3:0]    _zz_updatedEntry_3_srcReady_1_6;
  reg                 _zz_issueEntry_valid_4;
  reg        [4:0]    _zz_issueEntry_robIdx;
  reg        [31:0]   _zz_issueEntry_branchInfo_predictPC;
  reg                 _zz_issueEntry_branchInfo_predictResult;
  reg                 _zz_issueEntry_exceptionInfo_exception;
  reg        [5:0]    _zz_issueEntry_exceptionInfo_eCode;
  reg        [0:0]    _zz_issueEntry_exceptionInfo_eSubCode;
  reg        [31:0]   _zz_issueEntry_pc;
  reg        [5:0]    _zz_issueEntry_prd;
  reg        [5:0]    _zz_issueEntry_psrc_0;
  reg        [5:0]    _zz_issueEntry_psrc_1;
  reg        [31:0]   _zz_issueEntry_imm;
  reg        [3:0]    _zz_issueEntry_uop_aluOp;
  reg        [1:0]    _zz_issueEntry_uop_bruOp;
  reg        [1:0]    _zz_issueEntry_uop_cruOp;
  reg        [2:0]    _zz_issueEntry_roop_aluROOp;
  reg                 _zz_issueEntry_srcReady_0;
  reg                 _zz_issueEntry_srcReady_1;
  reg                 queue_0_valid;
  reg        [4:0]    queue_0_robIdx;
  reg        [31:0]   queue_0_branchInfo_predictPC;
  reg                 queue_0_branchInfo_predictResult;
  reg                 queue_0_exceptionInfo_exception;
  reg        [5:0]    queue_0_exceptionInfo_eCode;
  reg        [0:0]    queue_0_exceptionInfo_eSubCode;
  reg        [31:0]   queue_0_pc;
  reg        [5:0]    queue_0_prd;
  reg        [5:0]    queue_0_psrc_0;
  reg        [5:0]    queue_0_psrc_1;
  reg        [31:0]   queue_0_imm;
  reg        [3:0]    queue_0_uop_aluOp;
  reg        [1:0]    queue_0_uop_bruOp;
  reg        [1:0]    queue_0_uop_cruOp;
  reg        [2:0]    queue_0_roop_aluROOp;
  reg                 queue_0_srcReady_0;
  reg                 queue_0_srcReady_1;
  reg                 queue_1_valid;
  reg        [4:0]    queue_1_robIdx;
  reg        [31:0]   queue_1_branchInfo_predictPC;
  reg                 queue_1_branchInfo_predictResult;
  reg                 queue_1_exceptionInfo_exception;
  reg        [5:0]    queue_1_exceptionInfo_eCode;
  reg        [0:0]    queue_1_exceptionInfo_eSubCode;
  reg        [31:0]   queue_1_pc;
  reg        [5:0]    queue_1_prd;
  reg        [5:0]    queue_1_psrc_0;
  reg        [5:0]    queue_1_psrc_1;
  reg        [31:0]   queue_1_imm;
  reg        [3:0]    queue_1_uop_aluOp;
  reg        [1:0]    queue_1_uop_bruOp;
  reg        [1:0]    queue_1_uop_cruOp;
  reg        [2:0]    queue_1_roop_aluROOp;
  reg                 queue_1_srcReady_0;
  reg                 queue_1_srcReady_1;
  reg                 queue_2_valid;
  reg        [4:0]    queue_2_robIdx;
  reg        [31:0]   queue_2_branchInfo_predictPC;
  reg                 queue_2_branchInfo_predictResult;
  reg                 queue_2_exceptionInfo_exception;
  reg        [5:0]    queue_2_exceptionInfo_eCode;
  reg        [0:0]    queue_2_exceptionInfo_eSubCode;
  reg        [31:0]   queue_2_pc;
  reg        [5:0]    queue_2_prd;
  reg        [5:0]    queue_2_psrc_0;
  reg        [5:0]    queue_2_psrc_1;
  reg        [31:0]   queue_2_imm;
  reg        [3:0]    queue_2_uop_aluOp;
  reg        [1:0]    queue_2_uop_bruOp;
  reg        [1:0]    queue_2_uop_cruOp;
  reg        [2:0]    queue_2_roop_aluROOp;
  reg                 queue_2_srcReady_0;
  reg                 queue_2_srcReady_1;
  reg                 queue_3_valid;
  reg        [4:0]    queue_3_robIdx;
  reg        [31:0]   queue_3_branchInfo_predictPC;
  reg                 queue_3_branchInfo_predictResult;
  reg                 queue_3_exceptionInfo_exception;
  reg        [5:0]    queue_3_exceptionInfo_eCode;
  reg        [0:0]    queue_3_exceptionInfo_eSubCode;
  reg        [31:0]   queue_3_pc;
  reg        [5:0]    queue_3_prd;
  reg        [5:0]    queue_3_psrc_0;
  reg        [5:0]    queue_3_psrc_1;
  reg        [31:0]   queue_3_imm;
  reg        [3:0]    queue_3_uop_aluOp;
  reg        [1:0]    queue_3_uop_bruOp;
  reg        [1:0]    queue_3_uop_cruOp;
  reg        [2:0]    queue_3_roop_aluROOp;
  reg                 queue_3_srcReady_0;
  reg                 queue_3_srcReady_1;
  reg        [3:0]    readyToIssue;
  wire       [3:0]    readyToIssue_ohFirst_input;
  wire       [3:0]    readyToIssue_ohFirst_masked;
  wire       [3:0]    issueVector;
  reg        [3:0]    shiftAhead;
  reg        [4:0]    emptyEntry;
  wire       [4:0]    emptyEntry_ohFirst_input;
  wire       [4:0]    emptyEntry_ohFirst_masked;
  wire       [4:0]    writeVector;
  wire                updatedEntry_0_valid;
  wire       [4:0]    updatedEntry_0_robIdx;
  wire       [31:0]   updatedEntry_0_branchInfo_predictPC;
  wire                updatedEntry_0_branchInfo_predictResult;
  wire                updatedEntry_0_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_0_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_0_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_0_pc;
  wire       [5:0]    updatedEntry_0_prd;
  wire       [5:0]    updatedEntry_0_psrc_0;
  wire       [5:0]    updatedEntry_0_psrc_1;
  wire       [31:0]   updatedEntry_0_imm;
  wire       [3:0]    updatedEntry_0_uop_aluOp;
  wire       [1:0]    updatedEntry_0_uop_bruOp;
  wire       [1:0]    updatedEntry_0_uop_cruOp;
  wire       [2:0]    updatedEntry_0_roop_aluROOp;
  reg                 updatedEntry_0_srcReady_0;
  reg                 updatedEntry_0_srcReady_1;
  wire                updatedEntry_1_valid;
  wire       [4:0]    updatedEntry_1_robIdx;
  wire       [31:0]   updatedEntry_1_branchInfo_predictPC;
  wire                updatedEntry_1_branchInfo_predictResult;
  wire                updatedEntry_1_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_1_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_1_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_1_pc;
  wire       [5:0]    updatedEntry_1_prd;
  wire       [5:0]    updatedEntry_1_psrc_0;
  wire       [5:0]    updatedEntry_1_psrc_1;
  wire       [31:0]   updatedEntry_1_imm;
  wire       [3:0]    updatedEntry_1_uop_aluOp;
  wire       [1:0]    updatedEntry_1_uop_bruOp;
  wire       [1:0]    updatedEntry_1_uop_cruOp;
  wire       [2:0]    updatedEntry_1_roop_aluROOp;
  reg                 updatedEntry_1_srcReady_0;
  reg                 updatedEntry_1_srcReady_1;
  wire                updatedEntry_2_valid;
  wire       [4:0]    updatedEntry_2_robIdx;
  wire       [31:0]   updatedEntry_2_branchInfo_predictPC;
  wire                updatedEntry_2_branchInfo_predictResult;
  wire                updatedEntry_2_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_2_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_2_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_2_pc;
  wire       [5:0]    updatedEntry_2_prd;
  wire       [5:0]    updatedEntry_2_psrc_0;
  wire       [5:0]    updatedEntry_2_psrc_1;
  wire       [31:0]   updatedEntry_2_imm;
  wire       [3:0]    updatedEntry_2_uop_aluOp;
  wire       [1:0]    updatedEntry_2_uop_bruOp;
  wire       [1:0]    updatedEntry_2_uop_cruOp;
  wire       [2:0]    updatedEntry_2_roop_aluROOp;
  reg                 updatedEntry_2_srcReady_0;
  reg                 updatedEntry_2_srcReady_1;
  wire                updatedEntry_3_valid;
  wire       [4:0]    updatedEntry_3_robIdx;
  wire       [31:0]   updatedEntry_3_branchInfo_predictPC;
  wire                updatedEntry_3_branchInfo_predictResult;
  wire                updatedEntry_3_exceptionInfo_exception;
  wire       [5:0]    updatedEntry_3_exceptionInfo_eCode;
  wire       [0:0]    updatedEntry_3_exceptionInfo_eSubCode;
  wire       [31:0]   updatedEntry_3_pc;
  wire       [5:0]    updatedEntry_3_prd;
  wire       [5:0]    updatedEntry_3_psrc_0;
  wire       [5:0]    updatedEntry_3_psrc_1;
  wire       [31:0]   updatedEntry_3_imm;
  wire       [3:0]    updatedEntry_3_uop_aluOp;
  wire       [1:0]    updatedEntry_3_uop_bruOp;
  wire       [1:0]    updatedEntry_3_uop_cruOp;
  wire       [2:0]    updatedEntry_3_roop_aluROOp;
  reg                 updatedEntry_3_srcReady_0;
  reg                 updatedEntry_3_srcReady_1;
  wire                appendEntry_valid;
  wire       [4:0]    appendEntry_robIdx;
  wire       [31:0]   appendEntry_branchInfo_predictPC;
  wire                appendEntry_branchInfo_predictResult;
  wire                appendEntry_exceptionInfo_exception;
  wire       [5:0]    appendEntry_exceptionInfo_eCode;
  wire       [0:0]    appendEntry_exceptionInfo_eSubCode;
  wire       [31:0]   appendEntry_pc;
  wire       [5:0]    appendEntry_prd;
  wire       [5:0]    appendEntry_psrc_0;
  wire       [5:0]    appendEntry_psrc_1;
  wire       [31:0]   appendEntry_imm;
  wire       [3:0]    appendEntry_uop_aluOp;
  wire       [1:0]    appendEntry_uop_bruOp;
  wire       [1:0]    appendEntry_uop_cruOp;
  wire       [2:0]    appendEntry_roop_aluROOp;
  wire                appendEntry_srcReady_0;
  wire                appendEntry_srcReady_1;
  reg                 queueNext_0_valid;
  reg        [4:0]    queueNext_0_robIdx;
  reg        [31:0]   queueNext_0_branchInfo_predictPC;
  reg                 queueNext_0_branchInfo_predictResult;
  reg                 queueNext_0_exceptionInfo_exception;
  reg        [5:0]    queueNext_0_exceptionInfo_eCode;
  reg        [0:0]    queueNext_0_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_0_pc;
  reg        [5:0]    queueNext_0_prd;
  reg        [5:0]    queueNext_0_psrc_0;
  reg        [5:0]    queueNext_0_psrc_1;
  reg        [31:0]   queueNext_0_imm;
  reg        [3:0]    queueNext_0_uop_aluOp;
  reg        [1:0]    queueNext_0_uop_bruOp;
  reg        [1:0]    queueNext_0_uop_cruOp;
  reg        [2:0]    queueNext_0_roop_aluROOp;
  reg                 queueNext_0_srcReady_0;
  reg                 queueNext_0_srcReady_1;
  reg                 queueNext_1_valid;
  reg        [4:0]    queueNext_1_robIdx;
  reg        [31:0]   queueNext_1_branchInfo_predictPC;
  reg                 queueNext_1_branchInfo_predictResult;
  reg                 queueNext_1_exceptionInfo_exception;
  reg        [5:0]    queueNext_1_exceptionInfo_eCode;
  reg        [0:0]    queueNext_1_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_1_pc;
  reg        [5:0]    queueNext_1_prd;
  reg        [5:0]    queueNext_1_psrc_0;
  reg        [5:0]    queueNext_1_psrc_1;
  reg        [31:0]   queueNext_1_imm;
  reg        [3:0]    queueNext_1_uop_aluOp;
  reg        [1:0]    queueNext_1_uop_bruOp;
  reg        [1:0]    queueNext_1_uop_cruOp;
  reg        [2:0]    queueNext_1_roop_aluROOp;
  reg                 queueNext_1_srcReady_0;
  reg                 queueNext_1_srcReady_1;
  reg                 queueNext_2_valid;
  reg        [4:0]    queueNext_2_robIdx;
  reg        [31:0]   queueNext_2_branchInfo_predictPC;
  reg                 queueNext_2_branchInfo_predictResult;
  reg                 queueNext_2_exceptionInfo_exception;
  reg        [5:0]    queueNext_2_exceptionInfo_eCode;
  reg        [0:0]    queueNext_2_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_2_pc;
  reg        [5:0]    queueNext_2_prd;
  reg        [5:0]    queueNext_2_psrc_0;
  reg        [5:0]    queueNext_2_psrc_1;
  reg        [31:0]   queueNext_2_imm;
  reg        [3:0]    queueNext_2_uop_aluOp;
  reg        [1:0]    queueNext_2_uop_bruOp;
  reg        [1:0]    queueNext_2_uop_cruOp;
  reg        [2:0]    queueNext_2_roop_aluROOp;
  reg                 queueNext_2_srcReady_0;
  reg                 queueNext_2_srcReady_1;
  reg                 queueNext_3_valid;
  reg        [4:0]    queueNext_3_robIdx;
  reg        [31:0]   queueNext_3_branchInfo_predictPC;
  reg                 queueNext_3_branchInfo_predictResult;
  reg                 queueNext_3_exceptionInfo_exception;
  reg        [5:0]    queueNext_3_exceptionInfo_eCode;
  reg        [0:0]    queueNext_3_exceptionInfo_eSubCode;
  reg        [31:0]   queueNext_3_pc;
  reg        [5:0]    queueNext_3_prd;
  reg        [5:0]    queueNext_3_psrc_0;
  reg        [5:0]    queueNext_3_psrc_1;
  reg        [31:0]   queueNext_3_imm;
  reg        [3:0]    queueNext_3_uop_aluOp;
  reg        [1:0]    queueNext_3_uop_bruOp;
  reg        [1:0]    queueNext_3_uop_cruOp;
  reg        [2:0]    queueNext_3_roop_aluROOp;
  reg                 queueNext_3_srcReady_0;
  reg                 queueNext_3_srcReady_1;
  wire                when_IssueQueue_l81;
  wire                when_IssueQueue_l83;
  wire                when_IssueQueue_l96;
  wire                when_IssueQueue_l81_1;
  wire                when_IssueQueue_l83_1;
  wire                when_IssueQueue_l96_1;
  wire                when_IssueQueue_l81_2;
  wire                when_IssueQueue_l83_2;
  wire                when_IssueQueue_l96_2;
  wire                when_IssueQueue_l81_3;
  wire                when_IssueQueue_l89;
  wire                when_IssueQueue_l96_3;
  reg        [3:0]    _zz_io_csrInQueue;
  wire                io_output_fire;
  wire                _zz_issueEntry_valid;
  wire                _zz_issueEntry_valid_1;
  wire                _zz_issueEntry_valid_2;
  wire       [1:0]    _zz_issueEntry_valid_3;
  wire                issueEntry_valid;
  wire       [4:0]    issueEntry_robIdx;
  wire       [31:0]   issueEntry_branchInfo_predictPC;
  wire                issueEntry_branchInfo_predictResult;
  wire                issueEntry_exceptionInfo_exception;
  wire       [5:0]    issueEntry_exceptionInfo_eCode;
  wire       [0:0]    issueEntry_exceptionInfo_eSubCode;
  wire       [31:0]   issueEntry_pc;
  wire       [5:0]    issueEntry_prd;
  wire       [5:0]    issueEntry_psrc_0;
  wire       [5:0]    issueEntry_psrc_1;
  wire       [31:0]   issueEntry_imm;
  wire       [3:0]    issueEntry_uop_aluOp;
  wire       [1:0]    issueEntry_uop_bruOp;
  wire       [1:0]    issueEntry_uop_cruOp;
  wire       [2:0]    issueEntry_roop_aluROOp;
  wire                issueEntry_srcReady_0;
  wire                issueEntry_srcReady_1;
  `ifndef SYNTHESIS
  reg [39:0] io_input_payload_uop_aluOp_string;
  reg [39:0] io_input_payload_uop_bruOp_string;
  reg [31:0] io_input_payload_uop_cruOp_string;
  reg [55:0] io_input_payload_roop_aluROOp_string;
  reg [39:0] io_output_payload_uop_aluOp_string;
  reg [39:0] io_output_payload_uop_bruOp_string;
  reg [31:0] io_output_payload_uop_cruOp_string;
  reg [55:0] io_output_payload_roop_aluROOp_string;
  reg [39:0] queue_0_uop_aluOp_string;
  reg [39:0] queue_0_uop_bruOp_string;
  reg [31:0] queue_0_uop_cruOp_string;
  reg [55:0] queue_0_roop_aluROOp_string;
  reg [39:0] queue_1_uop_aluOp_string;
  reg [39:0] queue_1_uop_bruOp_string;
  reg [31:0] queue_1_uop_cruOp_string;
  reg [55:0] queue_1_roop_aluROOp_string;
  reg [39:0] queue_2_uop_aluOp_string;
  reg [39:0] queue_2_uop_bruOp_string;
  reg [31:0] queue_2_uop_cruOp_string;
  reg [55:0] queue_2_roop_aluROOp_string;
  reg [39:0] queue_3_uop_aluOp_string;
  reg [39:0] queue_3_uop_bruOp_string;
  reg [31:0] queue_3_uop_cruOp_string;
  reg [55:0] queue_3_roop_aluROOp_string;
  reg [39:0] updatedEntry_0_uop_aluOp_string;
  reg [39:0] updatedEntry_0_uop_bruOp_string;
  reg [31:0] updatedEntry_0_uop_cruOp_string;
  reg [55:0] updatedEntry_0_roop_aluROOp_string;
  reg [39:0] updatedEntry_1_uop_aluOp_string;
  reg [39:0] updatedEntry_1_uop_bruOp_string;
  reg [31:0] updatedEntry_1_uop_cruOp_string;
  reg [55:0] updatedEntry_1_roop_aluROOp_string;
  reg [39:0] updatedEntry_2_uop_aluOp_string;
  reg [39:0] updatedEntry_2_uop_bruOp_string;
  reg [31:0] updatedEntry_2_uop_cruOp_string;
  reg [55:0] updatedEntry_2_roop_aluROOp_string;
  reg [39:0] updatedEntry_3_uop_aluOp_string;
  reg [39:0] updatedEntry_3_uop_bruOp_string;
  reg [31:0] updatedEntry_3_uop_cruOp_string;
  reg [55:0] updatedEntry_3_roop_aluROOp_string;
  reg [39:0] appendEntry_uop_aluOp_string;
  reg [39:0] appendEntry_uop_bruOp_string;
  reg [31:0] appendEntry_uop_cruOp_string;
  reg [55:0] appendEntry_roop_aluROOp_string;
  reg [39:0] queueNext_0_uop_aluOp_string;
  reg [39:0] queueNext_0_uop_bruOp_string;
  reg [31:0] queueNext_0_uop_cruOp_string;
  reg [55:0] queueNext_0_roop_aluROOp_string;
  reg [39:0] queueNext_1_uop_aluOp_string;
  reg [39:0] queueNext_1_uop_bruOp_string;
  reg [31:0] queueNext_1_uop_cruOp_string;
  reg [55:0] queueNext_1_roop_aluROOp_string;
  reg [39:0] queueNext_2_uop_aluOp_string;
  reg [39:0] queueNext_2_uop_bruOp_string;
  reg [31:0] queueNext_2_uop_cruOp_string;
  reg [55:0] queueNext_2_roop_aluROOp_string;
  reg [39:0] queueNext_3_uop_aluOp_string;
  reg [39:0] queueNext_3_uop_bruOp_string;
  reg [31:0] queueNext_3_uop_cruOp_string;
  reg [55:0] queueNext_3_roop_aluROOp_string;
  reg [39:0] issueEntry_uop_aluOp_string;
  reg [39:0] issueEntry_uop_bruOp_string;
  reg [31:0] issueEntry_uop_cruOp_string;
  reg [55:0] issueEntry_roop_aluROOp_string;
  `endif


  assign _zz_readyToIssue_ohFirst_masked = (readyToIssue_ohFirst_input - 4'b0001);
  assign _zz_emptyEntry_ohFirst_masked = (emptyEntry_ohFirst_input - 5'h01);
  assign _zz_appendEntry_srcReady_0 = (io_input_payload_psrc_0 == io_writebackSignal_3);
  assign _zz_appendEntry_srcReady_0_1 = (io_input_payload_psrc_0 == io_writebackSignal_2);
  assign _zz_appendEntry_srcReady_0_2 = {(io_input_payload_psrc_0 == io_writebackSignal_1),(io_input_payload_psrc_0 == io_writebackSignal_0)};
  assign _zz_appendEntry_srcReady_0_3 = (io_input_payload_psrc_0 == io_earlyWakeup_7_payload);
  assign _zz_appendEntry_srcReady_0_4 = ((io_input_payload_psrc_0 == io_earlyWakeup_6_payload) && io_earlyWakeup_6_valid);
  assign _zz_appendEntry_srcReady_0_5 = ((io_input_payload_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_appendEntry_srcReady_0_6 = {((io_input_payload_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid),{(_zz_appendEntry_srcReady_0_7 && io_earlyWakeup_3_valid),{_zz_appendEntry_srcReady_0_8,{_zz_appendEntry_srcReady_0_9,_zz_appendEntry_srcReady_0_10}}}};
  assign _zz_appendEntry_srcReady_0_7 = (io_input_payload_psrc_0 == io_earlyWakeup_3_payload);
  assign _zz_appendEntry_srcReady_0_8 = ((io_input_payload_psrc_0 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid);
  assign _zz_appendEntry_srcReady_0_9 = ((io_input_payload_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid);
  assign _zz_appendEntry_srcReady_0_10 = ((io_input_payload_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid);
  assign _zz_appendEntry_srcReady_1 = (io_input_payload_psrc_1 == io_writebackSignal_2);
  assign _zz_appendEntry_srcReady_1_1 = (io_input_payload_psrc_1 == io_writebackSignal_1);
  assign _zz_appendEntry_srcReady_1_2 = (io_input_payload_psrc_1 == io_writebackSignal_0);
  assign _zz_appendEntry_srcReady_1_3 = (io_input_payload_psrc_1 == io_earlyWakeup_6_payload);
  assign _zz_appendEntry_srcReady_1_4 = ((io_input_payload_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_appendEntry_srcReady_1_5 = ((io_input_payload_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_appendEntry_srcReady_1_6 = {((io_input_payload_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((io_input_payload_psrc_1 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((io_input_payload_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((io_input_payload_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_0_srcReady_0 = (queue_0_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_0_srcReady_0_1 = (queue_0_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_0_srcReady_0_2 = (queue_0_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_0_srcReady_0_3 = (queue_0_psrc_0 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_0_srcReady_0_4 = ((queue_0_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_0_srcReady_0_5 = ((queue_0_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_0_srcReady_0_6 = {((queue_0_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_0_psrc_0 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_0_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_0_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_0_srcReady_1 = (queue_0_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_0_srcReady_1_1 = (queue_0_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_0_srcReady_1_2 = (queue_0_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_0_srcReady_1_3 = (queue_0_psrc_1 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_0_srcReady_1_4 = ((queue_0_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_0_srcReady_1_5 = ((queue_0_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_0_srcReady_1_6 = {((queue_0_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_0_psrc_1 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_0_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_0_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_1_srcReady_0 = (queue_1_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_1_srcReady_0_1 = (queue_1_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_1_srcReady_0_2 = (queue_1_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_1_srcReady_0_3 = (queue_1_psrc_0 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_1_srcReady_0_4 = ((queue_1_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_1_srcReady_0_5 = ((queue_1_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_1_srcReady_0_6 = {((queue_1_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_1_psrc_0 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_1_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_1_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_1_srcReady_1 = (queue_1_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_1_srcReady_1_1 = (queue_1_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_1_srcReady_1_2 = (queue_1_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_1_srcReady_1_3 = (queue_1_psrc_1 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_1_srcReady_1_4 = ((queue_1_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_1_srcReady_1_5 = ((queue_1_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_1_srcReady_1_6 = {((queue_1_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_1_psrc_1 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_1_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_1_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_2_srcReady_0 = (queue_2_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_2_srcReady_0_1 = (queue_2_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_2_srcReady_0_2 = (queue_2_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_2_srcReady_0_3 = (queue_2_psrc_0 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_2_srcReady_0_4 = ((queue_2_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_2_srcReady_0_5 = ((queue_2_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_2_srcReady_0_6 = {((queue_2_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_2_psrc_0 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_2_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_2_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_2_srcReady_1 = (queue_2_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_2_srcReady_1_1 = (queue_2_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_2_srcReady_1_2 = (queue_2_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_2_srcReady_1_3 = (queue_2_psrc_1 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_2_srcReady_1_4 = ((queue_2_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_2_srcReady_1_5 = ((queue_2_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_2_srcReady_1_6 = {((queue_2_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_2_psrc_1 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_2_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_2_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_3_srcReady_0 = (queue_3_psrc_0 == io_writebackSignal_2);
  assign _zz_updatedEntry_3_srcReady_0_1 = (queue_3_psrc_0 == io_writebackSignal_1);
  assign _zz_updatedEntry_3_srcReady_0_2 = (queue_3_psrc_0 == io_writebackSignal_0);
  assign _zz_updatedEntry_3_srcReady_0_3 = (queue_3_psrc_0 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_3_srcReady_0_4 = ((queue_3_psrc_0 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_3_srcReady_0_5 = ((queue_3_psrc_0 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_3_srcReady_0_6 = {((queue_3_psrc_0 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_3_psrc_0 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_3_psrc_0 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_3_psrc_0 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  assign _zz_updatedEntry_3_srcReady_1 = (queue_3_psrc_1 == io_writebackSignal_2);
  assign _zz_updatedEntry_3_srcReady_1_1 = (queue_3_psrc_1 == io_writebackSignal_1);
  assign _zz_updatedEntry_3_srcReady_1_2 = (queue_3_psrc_1 == io_writebackSignal_0);
  assign _zz_updatedEntry_3_srcReady_1_3 = (queue_3_psrc_1 == io_earlyWakeup_6_payload);
  assign _zz_updatedEntry_3_srcReady_1_4 = ((queue_3_psrc_1 == io_earlyWakeup_5_payload) && io_earlyWakeup_5_valid);
  assign _zz_updatedEntry_3_srcReady_1_5 = ((queue_3_psrc_1 == io_earlyWakeup_4_payload) && io_earlyWakeup_4_valid);
  assign _zz_updatedEntry_3_srcReady_1_6 = {((queue_3_psrc_1 == io_earlyWakeup_3_payload) && io_earlyWakeup_3_valid),{((queue_3_psrc_1 == io_earlyWakeup_2_payload) && io_earlyWakeup_2_valid),{((queue_3_psrc_1 == io_earlyWakeup_1_payload) && io_earlyWakeup_1_valid),((queue_3_psrc_1 == io_earlyWakeup_0_payload) && io_earlyWakeup_0_valid)}}};
  always @(*) begin
    case(_zz_issueEntry_valid_3)
      2'b00 : begin
        _zz_issueEntry_valid_4 = queue_0_valid;
        _zz_issueEntry_robIdx = queue_0_robIdx;
        _zz_issueEntry_branchInfo_predictPC = queue_0_branchInfo_predictPC;
        _zz_issueEntry_branchInfo_predictResult = queue_0_branchInfo_predictResult;
        _zz_issueEntry_exceptionInfo_exception = queue_0_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_0_pc;
        _zz_issueEntry_prd = queue_0_prd;
        _zz_issueEntry_psrc_0 = queue_0_psrc_0;
        _zz_issueEntry_psrc_1 = queue_0_psrc_1;
        _zz_issueEntry_imm = queue_0_imm;
        _zz_issueEntry_uop_aluOp = queue_0_uop_aluOp;
        _zz_issueEntry_uop_bruOp = queue_0_uop_bruOp;
        _zz_issueEntry_uop_cruOp = queue_0_uop_cruOp;
        _zz_issueEntry_roop_aluROOp = queue_0_roop_aluROOp;
        _zz_issueEntry_srcReady_0 = queue_0_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_0_srcReady_1;
      end
      2'b01 : begin
        _zz_issueEntry_valid_4 = queue_1_valid;
        _zz_issueEntry_robIdx = queue_1_robIdx;
        _zz_issueEntry_branchInfo_predictPC = queue_1_branchInfo_predictPC;
        _zz_issueEntry_branchInfo_predictResult = queue_1_branchInfo_predictResult;
        _zz_issueEntry_exceptionInfo_exception = queue_1_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_1_pc;
        _zz_issueEntry_prd = queue_1_prd;
        _zz_issueEntry_psrc_0 = queue_1_psrc_0;
        _zz_issueEntry_psrc_1 = queue_1_psrc_1;
        _zz_issueEntry_imm = queue_1_imm;
        _zz_issueEntry_uop_aluOp = queue_1_uop_aluOp;
        _zz_issueEntry_uop_bruOp = queue_1_uop_bruOp;
        _zz_issueEntry_uop_cruOp = queue_1_uop_cruOp;
        _zz_issueEntry_roop_aluROOp = queue_1_roop_aluROOp;
        _zz_issueEntry_srcReady_0 = queue_1_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_1_srcReady_1;
      end
      2'b10 : begin
        _zz_issueEntry_valid_4 = queue_2_valid;
        _zz_issueEntry_robIdx = queue_2_robIdx;
        _zz_issueEntry_branchInfo_predictPC = queue_2_branchInfo_predictPC;
        _zz_issueEntry_branchInfo_predictResult = queue_2_branchInfo_predictResult;
        _zz_issueEntry_exceptionInfo_exception = queue_2_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_2_pc;
        _zz_issueEntry_prd = queue_2_prd;
        _zz_issueEntry_psrc_0 = queue_2_psrc_0;
        _zz_issueEntry_psrc_1 = queue_2_psrc_1;
        _zz_issueEntry_imm = queue_2_imm;
        _zz_issueEntry_uop_aluOp = queue_2_uop_aluOp;
        _zz_issueEntry_uop_bruOp = queue_2_uop_bruOp;
        _zz_issueEntry_uop_cruOp = queue_2_uop_cruOp;
        _zz_issueEntry_roop_aluROOp = queue_2_roop_aluROOp;
        _zz_issueEntry_srcReady_0 = queue_2_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_2_srcReady_1;
      end
      default : begin
        _zz_issueEntry_valid_4 = queue_3_valid;
        _zz_issueEntry_robIdx = queue_3_robIdx;
        _zz_issueEntry_branchInfo_predictPC = queue_3_branchInfo_predictPC;
        _zz_issueEntry_branchInfo_predictResult = queue_3_branchInfo_predictResult;
        _zz_issueEntry_exceptionInfo_exception = queue_3_exceptionInfo_exception;
        _zz_issueEntry_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
        _zz_issueEntry_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
        _zz_issueEntry_pc = queue_3_pc;
        _zz_issueEntry_prd = queue_3_prd;
        _zz_issueEntry_psrc_0 = queue_3_psrc_0;
        _zz_issueEntry_psrc_1 = queue_3_psrc_1;
        _zz_issueEntry_imm = queue_3_imm;
        _zz_issueEntry_uop_aluOp = queue_3_uop_aluOp;
        _zz_issueEntry_uop_bruOp = queue_3_uop_bruOp;
        _zz_issueEntry_uop_cruOp = queue_3_uop_cruOp;
        _zz_issueEntry_roop_aluROOp = queue_3_roop_aluROOp;
        _zz_issueEntry_srcReady_0 = queue_3_srcReady_0;
        _zz_issueEntry_srcReady_1 = queue_3_srcReady_1;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_uop_aluOp)
      ALUOp_add : io_input_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_input_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_input_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_input_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_input_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_input_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_input_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_input_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_input_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_input_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_input_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_input_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_input_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_input_payload_uop_aluOp_string = "passb";
      default : io_input_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_input_payload_uop_bruOp)
      BRUOp_nop : io_input_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_input_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_input_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_input_payload_uop_bruOp_string = "ncadd";
      default : io_input_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_input_payload_uop_cruOp)
      CRUOp_nop : io_input_payload_uop_cruOp_string = "nop ";
      CRUOp_pass : io_input_payload_uop_cruOp_string = "pass";
      CRUOp_mask : io_input_payload_uop_cruOp_string = "mask";
      default : io_input_payload_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(io_input_payload_roop_aluROOp)
      ALUROOp_reg_1 : io_input_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : io_input_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : io_input_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : io_input_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : io_input_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : io_input_payload_roop_aluROOp_string = "linkreg";
      default : io_input_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_uop_aluOp)
      ALUOp_add : io_output_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_output_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_output_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_output_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_output_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_output_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_output_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_output_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_output_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_output_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_output_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_output_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_output_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_output_payload_uop_aluOp_string = "passb";
      default : io_output_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_uop_bruOp)
      BRUOp_nop : io_output_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_output_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_output_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_output_payload_uop_bruOp_string = "ncadd";
      default : io_output_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_uop_cruOp)
      CRUOp_nop : io_output_payload_uop_cruOp_string = "nop ";
      CRUOp_pass : io_output_payload_uop_cruOp_string = "pass";
      CRUOp_mask : io_output_payload_uop_cruOp_string = "mask";
      default : io_output_payload_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_roop_aluROOp)
      ALUROOp_reg_1 : io_output_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : io_output_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : io_output_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : io_output_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : io_output_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : io_output_payload_roop_aluROOp_string = "linkreg";
      default : io_output_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_0_uop_aluOp)
      ALUOp_add : queue_0_uop_aluOp_string = "add  ";
      ALUOp_sub : queue_0_uop_aluOp_string = "sub  ";
      ALUOp_slt : queue_0_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queue_0_uop_aluOp_string = "sltu ";
      ALUOp_eq : queue_0_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queue_0_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queue_0_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queue_0_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queue_0_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queue_0_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queue_0_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queue_0_uop_aluOp_string = "sra_1";
      ALUOp_passa : queue_0_uop_aluOp_string = "passa";
      ALUOp_passb : queue_0_uop_aluOp_string = "passb";
      default : queue_0_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_0_uop_bruOp)
      BRUOp_nop : queue_0_uop_bruOp_string = "nop  ";
      BRUOp_add : queue_0_uop_bruOp_string = "add  ";
      BRUOp_cadd : queue_0_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queue_0_uop_bruOp_string = "ncadd";
      default : queue_0_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_0_uop_cruOp)
      CRUOp_nop : queue_0_uop_cruOp_string = "nop ";
      CRUOp_pass : queue_0_uop_cruOp_string = "pass";
      CRUOp_mask : queue_0_uop_cruOp_string = "mask";
      default : queue_0_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(queue_0_roop_aluROOp)
      ALUROOp_reg_1 : queue_0_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queue_0_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queue_0_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queue_0_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queue_0_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queue_0_roop_aluROOp_string = "linkreg";
      default : queue_0_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_1_uop_aluOp)
      ALUOp_add : queue_1_uop_aluOp_string = "add  ";
      ALUOp_sub : queue_1_uop_aluOp_string = "sub  ";
      ALUOp_slt : queue_1_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queue_1_uop_aluOp_string = "sltu ";
      ALUOp_eq : queue_1_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queue_1_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queue_1_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queue_1_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queue_1_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queue_1_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queue_1_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queue_1_uop_aluOp_string = "sra_1";
      ALUOp_passa : queue_1_uop_aluOp_string = "passa";
      ALUOp_passb : queue_1_uop_aluOp_string = "passb";
      default : queue_1_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_1_uop_bruOp)
      BRUOp_nop : queue_1_uop_bruOp_string = "nop  ";
      BRUOp_add : queue_1_uop_bruOp_string = "add  ";
      BRUOp_cadd : queue_1_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queue_1_uop_bruOp_string = "ncadd";
      default : queue_1_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_1_uop_cruOp)
      CRUOp_nop : queue_1_uop_cruOp_string = "nop ";
      CRUOp_pass : queue_1_uop_cruOp_string = "pass";
      CRUOp_mask : queue_1_uop_cruOp_string = "mask";
      default : queue_1_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(queue_1_roop_aluROOp)
      ALUROOp_reg_1 : queue_1_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queue_1_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queue_1_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queue_1_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queue_1_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queue_1_roop_aluROOp_string = "linkreg";
      default : queue_1_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_2_uop_aluOp)
      ALUOp_add : queue_2_uop_aluOp_string = "add  ";
      ALUOp_sub : queue_2_uop_aluOp_string = "sub  ";
      ALUOp_slt : queue_2_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queue_2_uop_aluOp_string = "sltu ";
      ALUOp_eq : queue_2_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queue_2_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queue_2_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queue_2_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queue_2_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queue_2_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queue_2_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queue_2_uop_aluOp_string = "sra_1";
      ALUOp_passa : queue_2_uop_aluOp_string = "passa";
      ALUOp_passb : queue_2_uop_aluOp_string = "passb";
      default : queue_2_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_2_uop_bruOp)
      BRUOp_nop : queue_2_uop_bruOp_string = "nop  ";
      BRUOp_add : queue_2_uop_bruOp_string = "add  ";
      BRUOp_cadd : queue_2_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queue_2_uop_bruOp_string = "ncadd";
      default : queue_2_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_2_uop_cruOp)
      CRUOp_nop : queue_2_uop_cruOp_string = "nop ";
      CRUOp_pass : queue_2_uop_cruOp_string = "pass";
      CRUOp_mask : queue_2_uop_cruOp_string = "mask";
      default : queue_2_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(queue_2_roop_aluROOp)
      ALUROOp_reg_1 : queue_2_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queue_2_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queue_2_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queue_2_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queue_2_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queue_2_roop_aluROOp_string = "linkreg";
      default : queue_2_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queue_3_uop_aluOp)
      ALUOp_add : queue_3_uop_aluOp_string = "add  ";
      ALUOp_sub : queue_3_uop_aluOp_string = "sub  ";
      ALUOp_slt : queue_3_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queue_3_uop_aluOp_string = "sltu ";
      ALUOp_eq : queue_3_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queue_3_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queue_3_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queue_3_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queue_3_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queue_3_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queue_3_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queue_3_uop_aluOp_string = "sra_1";
      ALUOp_passa : queue_3_uop_aluOp_string = "passa";
      ALUOp_passb : queue_3_uop_aluOp_string = "passb";
      default : queue_3_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_3_uop_bruOp)
      BRUOp_nop : queue_3_uop_bruOp_string = "nop  ";
      BRUOp_add : queue_3_uop_bruOp_string = "add  ";
      BRUOp_cadd : queue_3_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queue_3_uop_bruOp_string = "ncadd";
      default : queue_3_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queue_3_uop_cruOp)
      CRUOp_nop : queue_3_uop_cruOp_string = "nop ";
      CRUOp_pass : queue_3_uop_cruOp_string = "pass";
      CRUOp_mask : queue_3_uop_cruOp_string = "mask";
      default : queue_3_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(queue_3_roop_aluROOp)
      ALUROOp_reg_1 : queue_3_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queue_3_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queue_3_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queue_3_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queue_3_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queue_3_roop_aluROOp_string = "linkreg";
      default : queue_3_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_uop_aluOp)
      ALUOp_add : updatedEntry_0_uop_aluOp_string = "add  ";
      ALUOp_sub : updatedEntry_0_uop_aluOp_string = "sub  ";
      ALUOp_slt : updatedEntry_0_uop_aluOp_string = "slt  ";
      ALUOp_sltu : updatedEntry_0_uop_aluOp_string = "sltu ";
      ALUOp_eq : updatedEntry_0_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : updatedEntry_0_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : updatedEntry_0_uop_aluOp_string = "and_1";
      ALUOp_or_1 : updatedEntry_0_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : updatedEntry_0_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : updatedEntry_0_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : updatedEntry_0_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : updatedEntry_0_uop_aluOp_string = "sra_1";
      ALUOp_passa : updatedEntry_0_uop_aluOp_string = "passa";
      ALUOp_passb : updatedEntry_0_uop_aluOp_string = "passb";
      default : updatedEntry_0_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_uop_bruOp)
      BRUOp_nop : updatedEntry_0_uop_bruOp_string = "nop  ";
      BRUOp_add : updatedEntry_0_uop_bruOp_string = "add  ";
      BRUOp_cadd : updatedEntry_0_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : updatedEntry_0_uop_bruOp_string = "ncadd";
      default : updatedEntry_0_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_uop_cruOp)
      CRUOp_nop : updatedEntry_0_uop_cruOp_string = "nop ";
      CRUOp_pass : updatedEntry_0_uop_cruOp_string = "pass";
      CRUOp_mask : updatedEntry_0_uop_cruOp_string = "mask";
      default : updatedEntry_0_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_0_roop_aluROOp)
      ALUROOp_reg_1 : updatedEntry_0_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : updatedEntry_0_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : updatedEntry_0_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : updatedEntry_0_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : updatedEntry_0_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : updatedEntry_0_roop_aluROOp_string = "linkreg";
      default : updatedEntry_0_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_uop_aluOp)
      ALUOp_add : updatedEntry_1_uop_aluOp_string = "add  ";
      ALUOp_sub : updatedEntry_1_uop_aluOp_string = "sub  ";
      ALUOp_slt : updatedEntry_1_uop_aluOp_string = "slt  ";
      ALUOp_sltu : updatedEntry_1_uop_aluOp_string = "sltu ";
      ALUOp_eq : updatedEntry_1_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : updatedEntry_1_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : updatedEntry_1_uop_aluOp_string = "and_1";
      ALUOp_or_1 : updatedEntry_1_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : updatedEntry_1_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : updatedEntry_1_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : updatedEntry_1_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : updatedEntry_1_uop_aluOp_string = "sra_1";
      ALUOp_passa : updatedEntry_1_uop_aluOp_string = "passa";
      ALUOp_passb : updatedEntry_1_uop_aluOp_string = "passb";
      default : updatedEntry_1_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_uop_bruOp)
      BRUOp_nop : updatedEntry_1_uop_bruOp_string = "nop  ";
      BRUOp_add : updatedEntry_1_uop_bruOp_string = "add  ";
      BRUOp_cadd : updatedEntry_1_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : updatedEntry_1_uop_bruOp_string = "ncadd";
      default : updatedEntry_1_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_uop_cruOp)
      CRUOp_nop : updatedEntry_1_uop_cruOp_string = "nop ";
      CRUOp_pass : updatedEntry_1_uop_cruOp_string = "pass";
      CRUOp_mask : updatedEntry_1_uop_cruOp_string = "mask";
      default : updatedEntry_1_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_1_roop_aluROOp)
      ALUROOp_reg_1 : updatedEntry_1_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : updatedEntry_1_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : updatedEntry_1_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : updatedEntry_1_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : updatedEntry_1_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : updatedEntry_1_roop_aluROOp_string = "linkreg";
      default : updatedEntry_1_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_uop_aluOp)
      ALUOp_add : updatedEntry_2_uop_aluOp_string = "add  ";
      ALUOp_sub : updatedEntry_2_uop_aluOp_string = "sub  ";
      ALUOp_slt : updatedEntry_2_uop_aluOp_string = "slt  ";
      ALUOp_sltu : updatedEntry_2_uop_aluOp_string = "sltu ";
      ALUOp_eq : updatedEntry_2_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : updatedEntry_2_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : updatedEntry_2_uop_aluOp_string = "and_1";
      ALUOp_or_1 : updatedEntry_2_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : updatedEntry_2_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : updatedEntry_2_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : updatedEntry_2_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : updatedEntry_2_uop_aluOp_string = "sra_1";
      ALUOp_passa : updatedEntry_2_uop_aluOp_string = "passa";
      ALUOp_passb : updatedEntry_2_uop_aluOp_string = "passb";
      default : updatedEntry_2_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_uop_bruOp)
      BRUOp_nop : updatedEntry_2_uop_bruOp_string = "nop  ";
      BRUOp_add : updatedEntry_2_uop_bruOp_string = "add  ";
      BRUOp_cadd : updatedEntry_2_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : updatedEntry_2_uop_bruOp_string = "ncadd";
      default : updatedEntry_2_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_uop_cruOp)
      CRUOp_nop : updatedEntry_2_uop_cruOp_string = "nop ";
      CRUOp_pass : updatedEntry_2_uop_cruOp_string = "pass";
      CRUOp_mask : updatedEntry_2_uop_cruOp_string = "mask";
      default : updatedEntry_2_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_2_roop_aluROOp)
      ALUROOp_reg_1 : updatedEntry_2_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : updatedEntry_2_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : updatedEntry_2_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : updatedEntry_2_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : updatedEntry_2_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : updatedEntry_2_roop_aluROOp_string = "linkreg";
      default : updatedEntry_2_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_uop_aluOp)
      ALUOp_add : updatedEntry_3_uop_aluOp_string = "add  ";
      ALUOp_sub : updatedEntry_3_uop_aluOp_string = "sub  ";
      ALUOp_slt : updatedEntry_3_uop_aluOp_string = "slt  ";
      ALUOp_sltu : updatedEntry_3_uop_aluOp_string = "sltu ";
      ALUOp_eq : updatedEntry_3_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : updatedEntry_3_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : updatedEntry_3_uop_aluOp_string = "and_1";
      ALUOp_or_1 : updatedEntry_3_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : updatedEntry_3_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : updatedEntry_3_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : updatedEntry_3_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : updatedEntry_3_uop_aluOp_string = "sra_1";
      ALUOp_passa : updatedEntry_3_uop_aluOp_string = "passa";
      ALUOp_passb : updatedEntry_3_uop_aluOp_string = "passb";
      default : updatedEntry_3_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_uop_bruOp)
      BRUOp_nop : updatedEntry_3_uop_bruOp_string = "nop  ";
      BRUOp_add : updatedEntry_3_uop_bruOp_string = "add  ";
      BRUOp_cadd : updatedEntry_3_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : updatedEntry_3_uop_bruOp_string = "ncadd";
      default : updatedEntry_3_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_uop_cruOp)
      CRUOp_nop : updatedEntry_3_uop_cruOp_string = "nop ";
      CRUOp_pass : updatedEntry_3_uop_cruOp_string = "pass";
      CRUOp_mask : updatedEntry_3_uop_cruOp_string = "mask";
      default : updatedEntry_3_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(updatedEntry_3_roop_aluROOp)
      ALUROOp_reg_1 : updatedEntry_3_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : updatedEntry_3_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : updatedEntry_3_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : updatedEntry_3_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : updatedEntry_3_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : updatedEntry_3_roop_aluROOp_string = "linkreg";
      default : updatedEntry_3_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(appendEntry_uop_aluOp)
      ALUOp_add : appendEntry_uop_aluOp_string = "add  ";
      ALUOp_sub : appendEntry_uop_aluOp_string = "sub  ";
      ALUOp_slt : appendEntry_uop_aluOp_string = "slt  ";
      ALUOp_sltu : appendEntry_uop_aluOp_string = "sltu ";
      ALUOp_eq : appendEntry_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : appendEntry_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : appendEntry_uop_aluOp_string = "and_1";
      ALUOp_or_1 : appendEntry_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : appendEntry_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : appendEntry_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : appendEntry_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : appendEntry_uop_aluOp_string = "sra_1";
      ALUOp_passa : appendEntry_uop_aluOp_string = "passa";
      ALUOp_passb : appendEntry_uop_aluOp_string = "passb";
      default : appendEntry_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(appendEntry_uop_bruOp)
      BRUOp_nop : appendEntry_uop_bruOp_string = "nop  ";
      BRUOp_add : appendEntry_uop_bruOp_string = "add  ";
      BRUOp_cadd : appendEntry_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : appendEntry_uop_bruOp_string = "ncadd";
      default : appendEntry_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(appendEntry_uop_cruOp)
      CRUOp_nop : appendEntry_uop_cruOp_string = "nop ";
      CRUOp_pass : appendEntry_uop_cruOp_string = "pass";
      CRUOp_mask : appendEntry_uop_cruOp_string = "mask";
      default : appendEntry_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(appendEntry_roop_aluROOp)
      ALUROOp_reg_1 : appendEntry_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : appendEntry_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : appendEntry_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : appendEntry_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : appendEntry_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : appendEntry_roop_aluROOp_string = "linkreg";
      default : appendEntry_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_0_uop_aluOp)
      ALUOp_add : queueNext_0_uop_aluOp_string = "add  ";
      ALUOp_sub : queueNext_0_uop_aluOp_string = "sub  ";
      ALUOp_slt : queueNext_0_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queueNext_0_uop_aluOp_string = "sltu ";
      ALUOp_eq : queueNext_0_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queueNext_0_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queueNext_0_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queueNext_0_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queueNext_0_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queueNext_0_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queueNext_0_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queueNext_0_uop_aluOp_string = "sra_1";
      ALUOp_passa : queueNext_0_uop_aluOp_string = "passa";
      ALUOp_passb : queueNext_0_uop_aluOp_string = "passb";
      default : queueNext_0_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_0_uop_bruOp)
      BRUOp_nop : queueNext_0_uop_bruOp_string = "nop  ";
      BRUOp_add : queueNext_0_uop_bruOp_string = "add  ";
      BRUOp_cadd : queueNext_0_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queueNext_0_uop_bruOp_string = "ncadd";
      default : queueNext_0_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_0_uop_cruOp)
      CRUOp_nop : queueNext_0_uop_cruOp_string = "nop ";
      CRUOp_pass : queueNext_0_uop_cruOp_string = "pass";
      CRUOp_mask : queueNext_0_uop_cruOp_string = "mask";
      default : queueNext_0_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(queueNext_0_roop_aluROOp)
      ALUROOp_reg_1 : queueNext_0_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queueNext_0_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queueNext_0_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queueNext_0_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queueNext_0_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queueNext_0_roop_aluROOp_string = "linkreg";
      default : queueNext_0_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_1_uop_aluOp)
      ALUOp_add : queueNext_1_uop_aluOp_string = "add  ";
      ALUOp_sub : queueNext_1_uop_aluOp_string = "sub  ";
      ALUOp_slt : queueNext_1_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queueNext_1_uop_aluOp_string = "sltu ";
      ALUOp_eq : queueNext_1_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queueNext_1_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queueNext_1_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queueNext_1_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queueNext_1_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queueNext_1_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queueNext_1_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queueNext_1_uop_aluOp_string = "sra_1";
      ALUOp_passa : queueNext_1_uop_aluOp_string = "passa";
      ALUOp_passb : queueNext_1_uop_aluOp_string = "passb";
      default : queueNext_1_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_1_uop_bruOp)
      BRUOp_nop : queueNext_1_uop_bruOp_string = "nop  ";
      BRUOp_add : queueNext_1_uop_bruOp_string = "add  ";
      BRUOp_cadd : queueNext_1_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queueNext_1_uop_bruOp_string = "ncadd";
      default : queueNext_1_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_1_uop_cruOp)
      CRUOp_nop : queueNext_1_uop_cruOp_string = "nop ";
      CRUOp_pass : queueNext_1_uop_cruOp_string = "pass";
      CRUOp_mask : queueNext_1_uop_cruOp_string = "mask";
      default : queueNext_1_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(queueNext_1_roop_aluROOp)
      ALUROOp_reg_1 : queueNext_1_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queueNext_1_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queueNext_1_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queueNext_1_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queueNext_1_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queueNext_1_roop_aluROOp_string = "linkreg";
      default : queueNext_1_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_2_uop_aluOp)
      ALUOp_add : queueNext_2_uop_aluOp_string = "add  ";
      ALUOp_sub : queueNext_2_uop_aluOp_string = "sub  ";
      ALUOp_slt : queueNext_2_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queueNext_2_uop_aluOp_string = "sltu ";
      ALUOp_eq : queueNext_2_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queueNext_2_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queueNext_2_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queueNext_2_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queueNext_2_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queueNext_2_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queueNext_2_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queueNext_2_uop_aluOp_string = "sra_1";
      ALUOp_passa : queueNext_2_uop_aluOp_string = "passa";
      ALUOp_passb : queueNext_2_uop_aluOp_string = "passb";
      default : queueNext_2_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_2_uop_bruOp)
      BRUOp_nop : queueNext_2_uop_bruOp_string = "nop  ";
      BRUOp_add : queueNext_2_uop_bruOp_string = "add  ";
      BRUOp_cadd : queueNext_2_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queueNext_2_uop_bruOp_string = "ncadd";
      default : queueNext_2_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_2_uop_cruOp)
      CRUOp_nop : queueNext_2_uop_cruOp_string = "nop ";
      CRUOp_pass : queueNext_2_uop_cruOp_string = "pass";
      CRUOp_mask : queueNext_2_uop_cruOp_string = "mask";
      default : queueNext_2_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(queueNext_2_roop_aluROOp)
      ALUROOp_reg_1 : queueNext_2_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queueNext_2_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queueNext_2_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queueNext_2_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queueNext_2_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queueNext_2_roop_aluROOp_string = "linkreg";
      default : queueNext_2_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(queueNext_3_uop_aluOp)
      ALUOp_add : queueNext_3_uop_aluOp_string = "add  ";
      ALUOp_sub : queueNext_3_uop_aluOp_string = "sub  ";
      ALUOp_slt : queueNext_3_uop_aluOp_string = "slt  ";
      ALUOp_sltu : queueNext_3_uop_aluOp_string = "sltu ";
      ALUOp_eq : queueNext_3_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : queueNext_3_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : queueNext_3_uop_aluOp_string = "and_1";
      ALUOp_or_1 : queueNext_3_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : queueNext_3_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : queueNext_3_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : queueNext_3_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : queueNext_3_uop_aluOp_string = "sra_1";
      ALUOp_passa : queueNext_3_uop_aluOp_string = "passa";
      ALUOp_passb : queueNext_3_uop_aluOp_string = "passb";
      default : queueNext_3_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_3_uop_bruOp)
      BRUOp_nop : queueNext_3_uop_bruOp_string = "nop  ";
      BRUOp_add : queueNext_3_uop_bruOp_string = "add  ";
      BRUOp_cadd : queueNext_3_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : queueNext_3_uop_bruOp_string = "ncadd";
      default : queueNext_3_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(queueNext_3_uop_cruOp)
      CRUOp_nop : queueNext_3_uop_cruOp_string = "nop ";
      CRUOp_pass : queueNext_3_uop_cruOp_string = "pass";
      CRUOp_mask : queueNext_3_uop_cruOp_string = "mask";
      default : queueNext_3_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(queueNext_3_roop_aluROOp)
      ALUROOp_reg_1 : queueNext_3_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : queueNext_3_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : queueNext_3_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : queueNext_3_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : queueNext_3_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : queueNext_3_roop_aluROOp_string = "linkreg";
      default : queueNext_3_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(issueEntry_uop_aluOp)
      ALUOp_add : issueEntry_uop_aluOp_string = "add  ";
      ALUOp_sub : issueEntry_uop_aluOp_string = "sub  ";
      ALUOp_slt : issueEntry_uop_aluOp_string = "slt  ";
      ALUOp_sltu : issueEntry_uop_aluOp_string = "sltu ";
      ALUOp_eq : issueEntry_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : issueEntry_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : issueEntry_uop_aluOp_string = "and_1";
      ALUOp_or_1 : issueEntry_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : issueEntry_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : issueEntry_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : issueEntry_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : issueEntry_uop_aluOp_string = "sra_1";
      ALUOp_passa : issueEntry_uop_aluOp_string = "passa";
      ALUOp_passb : issueEntry_uop_aluOp_string = "passb";
      default : issueEntry_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(issueEntry_uop_bruOp)
      BRUOp_nop : issueEntry_uop_bruOp_string = "nop  ";
      BRUOp_add : issueEntry_uop_bruOp_string = "add  ";
      BRUOp_cadd : issueEntry_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : issueEntry_uop_bruOp_string = "ncadd";
      default : issueEntry_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(issueEntry_uop_cruOp)
      CRUOp_nop : issueEntry_uop_cruOp_string = "nop ";
      CRUOp_pass : issueEntry_uop_cruOp_string = "pass";
      CRUOp_mask : issueEntry_uop_cruOp_string = "mask";
      default : issueEntry_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(issueEntry_roop_aluROOp)
      ALUROOp_reg_1 : issueEntry_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : issueEntry_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : issueEntry_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : issueEntry_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : issueEntry_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : issueEntry_roop_aluROOp_string = "linkreg";
      default : issueEntry_roop_aluROOp_string = "???????";
    endcase
  end
  `endif

  always @(*) begin
    readyToIssue[0] = ((queue_0_valid && queue_0_srcReady_0) && queue_0_srcReady_1);
    readyToIssue[1] = ((queue_1_valid && queue_1_srcReady_0) && queue_1_srcReady_1);
    readyToIssue[2] = ((queue_2_valid && queue_2_srcReady_0) && queue_2_srcReady_1);
    readyToIssue[3] = ((queue_3_valid && queue_3_srcReady_0) && queue_3_srcReady_1);
  end

  assign readyToIssue_ohFirst_input = readyToIssue;
  assign readyToIssue_ohFirst_masked = (readyToIssue_ohFirst_input & (~ _zz_readyToIssue_ohFirst_masked));
  assign issueVector = readyToIssue_ohFirst_masked;
  always @(*) begin
    emptyEntry[0] = (! queue_0_valid);
    emptyEntry[1] = (! queue_1_valid);
    emptyEntry[2] = (! queue_2_valid);
    emptyEntry[3] = (! queue_3_valid);
    emptyEntry[4] = 1'b1;
    emptyEntry[0] = (! queue_0_valid);
    emptyEntry[1] = (! queue_1_valid);
    emptyEntry[2] = (! queue_2_valid);
    emptyEntry[3] = (! queue_3_valid);
  end

  assign emptyEntry_ohFirst_input = emptyEntry;
  assign emptyEntry_ohFirst_masked = (emptyEntry_ohFirst_input & (~ _zz_emptyEntry_ohFirst_masked));
  assign writeVector = emptyEntry_ohFirst_masked;
  assign appendEntry_valid = io_input_valid;
  assign appendEntry_robIdx = io_input_payload_robIdx;
  assign appendEntry_branchInfo_predictPC = io_input_payload_branchInfo_predictPC;
  assign appendEntry_branchInfo_predictResult = io_input_payload_branchInfo_predictResult;
  assign appendEntry_exceptionInfo_exception = io_input_payload_exceptionInfo_exception;
  assign appendEntry_exceptionInfo_eCode = io_input_payload_exceptionInfo_eCode;
  assign appendEntry_exceptionInfo_eSubCode = io_input_payload_exceptionInfo_eSubCode;
  assign appendEntry_pc = io_input_payload_pc;
  assign appendEntry_prd = io_input_payload_prd;
  assign appendEntry_psrc_0 = io_input_payload_psrc_0;
  assign appendEntry_psrc_1 = io_input_payload_psrc_1;
  assign appendEntry_imm = io_input_payload_imm;
  assign appendEntry_uop_aluOp = io_input_payload_uop_aluOp;
  assign appendEntry_uop_bruOp = io_input_payload_uop_bruOp;
  assign appendEntry_uop_cruOp = io_input_payload_uop_cruOp;
  assign appendEntry_roop_aluROOp = io_input_payload_roop_aluROOp;
  assign appendEntry_srcReady_0 = ((io_input_payload_srcReady_0 || (|{(io_input_payload_psrc_0 == io_writebackSignal_4),{_zz_appendEntry_srcReady_0,{_zz_appendEntry_srcReady_0_1,_zz_appendEntry_srcReady_0_2}}})) || ((|{(_zz_appendEntry_srcReady_0_3 && io_earlyWakeup_7_valid),{_zz_appendEntry_srcReady_0_4,{_zz_appendEntry_srcReady_0_5,_zz_appendEntry_srcReady_0_6}}}) || ((io_input_payload_psrc_0 == io_wakeOut_payload) && io_wakeOut_valid)));
  assign appendEntry_srcReady_1 = ((io_input_payload_srcReady_1 || (|{(io_input_payload_psrc_1 == io_writebackSignal_4),{(io_input_payload_psrc_1 == io_writebackSignal_3),{_zz_appendEntry_srcReady_1,{_zz_appendEntry_srcReady_1_1,_zz_appendEntry_srcReady_1_2}}}})) || ((|{((io_input_payload_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_appendEntry_srcReady_1_3 && io_earlyWakeup_6_valid),{_zz_appendEntry_srcReady_1_4,{_zz_appendEntry_srcReady_1_5,_zz_appendEntry_srcReady_1_6}}}}) || ((io_input_payload_psrc_1 == io_wakeOut_payload) && io_wakeOut_valid)));
  assign updatedEntry_0_valid = queue_0_valid;
  assign updatedEntry_0_robIdx = queue_0_robIdx;
  assign updatedEntry_0_branchInfo_predictPC = queue_0_branchInfo_predictPC;
  assign updatedEntry_0_branchInfo_predictResult = queue_0_branchInfo_predictResult;
  assign updatedEntry_0_exceptionInfo_exception = queue_0_exceptionInfo_exception;
  assign updatedEntry_0_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
  assign updatedEntry_0_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
  assign updatedEntry_0_pc = queue_0_pc;
  assign updatedEntry_0_prd = queue_0_prd;
  assign updatedEntry_0_psrc_0 = queue_0_psrc_0;
  assign updatedEntry_0_psrc_1 = queue_0_psrc_1;
  assign updatedEntry_0_imm = queue_0_imm;
  assign updatedEntry_0_uop_aluOp = queue_0_uop_aluOp;
  assign updatedEntry_0_uop_bruOp = queue_0_uop_bruOp;
  assign updatedEntry_0_uop_cruOp = queue_0_uop_cruOp;
  assign updatedEntry_0_roop_aluROOp = queue_0_roop_aluROOp;
  always @(*) begin
    updatedEntry_0_srcReady_0 = queue_0_srcReady_0;
    updatedEntry_0_srcReady_0 = ((queue_0_srcReady_0 || (|{(queue_0_psrc_0 == io_writebackSignal_4),{(queue_0_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_0_srcReady_0,{_zz_updatedEntry_0_srcReady_0_1,_zz_updatedEntry_0_srcReady_0_2}}}})) || ((|{((queue_0_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_0_srcReady_0_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_0_srcReady_0_4,{_zz_updatedEntry_0_srcReady_0_5,_zz_updatedEntry_0_srcReady_0_6}}}}) || ((queue_0_psrc_0 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  always @(*) begin
    updatedEntry_0_srcReady_1 = queue_0_srcReady_1;
    updatedEntry_0_srcReady_1 = ((queue_0_srcReady_1 || (|{(queue_0_psrc_1 == io_writebackSignal_4),{(queue_0_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_0_srcReady_1,{_zz_updatedEntry_0_srcReady_1_1,_zz_updatedEntry_0_srcReady_1_2}}}})) || ((|{((queue_0_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_0_srcReady_1_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_0_srcReady_1_4,{_zz_updatedEntry_0_srcReady_1_5,_zz_updatedEntry_0_srcReady_1_6}}}}) || ((queue_0_psrc_1 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  assign updatedEntry_1_valid = queue_1_valid;
  assign updatedEntry_1_robIdx = queue_1_robIdx;
  assign updatedEntry_1_branchInfo_predictPC = queue_1_branchInfo_predictPC;
  assign updatedEntry_1_branchInfo_predictResult = queue_1_branchInfo_predictResult;
  assign updatedEntry_1_exceptionInfo_exception = queue_1_exceptionInfo_exception;
  assign updatedEntry_1_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
  assign updatedEntry_1_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
  assign updatedEntry_1_pc = queue_1_pc;
  assign updatedEntry_1_prd = queue_1_prd;
  assign updatedEntry_1_psrc_0 = queue_1_psrc_0;
  assign updatedEntry_1_psrc_1 = queue_1_psrc_1;
  assign updatedEntry_1_imm = queue_1_imm;
  assign updatedEntry_1_uop_aluOp = queue_1_uop_aluOp;
  assign updatedEntry_1_uop_bruOp = queue_1_uop_bruOp;
  assign updatedEntry_1_uop_cruOp = queue_1_uop_cruOp;
  assign updatedEntry_1_roop_aluROOp = queue_1_roop_aluROOp;
  always @(*) begin
    updatedEntry_1_srcReady_0 = queue_1_srcReady_0;
    updatedEntry_1_srcReady_0 = ((queue_1_srcReady_0 || (|{(queue_1_psrc_0 == io_writebackSignal_4),{(queue_1_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_1_srcReady_0,{_zz_updatedEntry_1_srcReady_0_1,_zz_updatedEntry_1_srcReady_0_2}}}})) || ((|{((queue_1_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_1_srcReady_0_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_1_srcReady_0_4,{_zz_updatedEntry_1_srcReady_0_5,_zz_updatedEntry_1_srcReady_0_6}}}}) || ((queue_1_psrc_0 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  always @(*) begin
    updatedEntry_1_srcReady_1 = queue_1_srcReady_1;
    updatedEntry_1_srcReady_1 = ((queue_1_srcReady_1 || (|{(queue_1_psrc_1 == io_writebackSignal_4),{(queue_1_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_1_srcReady_1,{_zz_updatedEntry_1_srcReady_1_1,_zz_updatedEntry_1_srcReady_1_2}}}})) || ((|{((queue_1_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_1_srcReady_1_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_1_srcReady_1_4,{_zz_updatedEntry_1_srcReady_1_5,_zz_updatedEntry_1_srcReady_1_6}}}}) || ((queue_1_psrc_1 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  assign updatedEntry_2_valid = queue_2_valid;
  assign updatedEntry_2_robIdx = queue_2_robIdx;
  assign updatedEntry_2_branchInfo_predictPC = queue_2_branchInfo_predictPC;
  assign updatedEntry_2_branchInfo_predictResult = queue_2_branchInfo_predictResult;
  assign updatedEntry_2_exceptionInfo_exception = queue_2_exceptionInfo_exception;
  assign updatedEntry_2_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
  assign updatedEntry_2_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
  assign updatedEntry_2_pc = queue_2_pc;
  assign updatedEntry_2_prd = queue_2_prd;
  assign updatedEntry_2_psrc_0 = queue_2_psrc_0;
  assign updatedEntry_2_psrc_1 = queue_2_psrc_1;
  assign updatedEntry_2_imm = queue_2_imm;
  assign updatedEntry_2_uop_aluOp = queue_2_uop_aluOp;
  assign updatedEntry_2_uop_bruOp = queue_2_uop_bruOp;
  assign updatedEntry_2_uop_cruOp = queue_2_uop_cruOp;
  assign updatedEntry_2_roop_aluROOp = queue_2_roop_aluROOp;
  always @(*) begin
    updatedEntry_2_srcReady_0 = queue_2_srcReady_0;
    updatedEntry_2_srcReady_0 = ((queue_2_srcReady_0 || (|{(queue_2_psrc_0 == io_writebackSignal_4),{(queue_2_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_2_srcReady_0,{_zz_updatedEntry_2_srcReady_0_1,_zz_updatedEntry_2_srcReady_0_2}}}})) || ((|{((queue_2_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_2_srcReady_0_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_2_srcReady_0_4,{_zz_updatedEntry_2_srcReady_0_5,_zz_updatedEntry_2_srcReady_0_6}}}}) || ((queue_2_psrc_0 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  always @(*) begin
    updatedEntry_2_srcReady_1 = queue_2_srcReady_1;
    updatedEntry_2_srcReady_1 = ((queue_2_srcReady_1 || (|{(queue_2_psrc_1 == io_writebackSignal_4),{(queue_2_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_2_srcReady_1,{_zz_updatedEntry_2_srcReady_1_1,_zz_updatedEntry_2_srcReady_1_2}}}})) || ((|{((queue_2_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_2_srcReady_1_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_2_srcReady_1_4,{_zz_updatedEntry_2_srcReady_1_5,_zz_updatedEntry_2_srcReady_1_6}}}}) || ((queue_2_psrc_1 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  assign updatedEntry_3_valid = queue_3_valid;
  assign updatedEntry_3_robIdx = queue_3_robIdx;
  assign updatedEntry_3_branchInfo_predictPC = queue_3_branchInfo_predictPC;
  assign updatedEntry_3_branchInfo_predictResult = queue_3_branchInfo_predictResult;
  assign updatedEntry_3_exceptionInfo_exception = queue_3_exceptionInfo_exception;
  assign updatedEntry_3_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
  assign updatedEntry_3_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
  assign updatedEntry_3_pc = queue_3_pc;
  assign updatedEntry_3_prd = queue_3_prd;
  assign updatedEntry_3_psrc_0 = queue_3_psrc_0;
  assign updatedEntry_3_psrc_1 = queue_3_psrc_1;
  assign updatedEntry_3_imm = queue_3_imm;
  assign updatedEntry_3_uop_aluOp = queue_3_uop_aluOp;
  assign updatedEntry_3_uop_bruOp = queue_3_uop_bruOp;
  assign updatedEntry_3_uop_cruOp = queue_3_uop_cruOp;
  assign updatedEntry_3_roop_aluROOp = queue_3_roop_aluROOp;
  always @(*) begin
    updatedEntry_3_srcReady_0 = queue_3_srcReady_0;
    updatedEntry_3_srcReady_0 = ((queue_3_srcReady_0 || (|{(queue_3_psrc_0 == io_writebackSignal_4),{(queue_3_psrc_0 == io_writebackSignal_3),{_zz_updatedEntry_3_srcReady_0,{_zz_updatedEntry_3_srcReady_0_1,_zz_updatedEntry_3_srcReady_0_2}}}})) || ((|{((queue_3_psrc_0 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_3_srcReady_0_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_3_srcReady_0_4,{_zz_updatedEntry_3_srcReady_0_5,_zz_updatedEntry_3_srcReady_0_6}}}}) || ((queue_3_psrc_0 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  always @(*) begin
    updatedEntry_3_srcReady_1 = queue_3_srcReady_1;
    updatedEntry_3_srcReady_1 = ((queue_3_srcReady_1 || (|{(queue_3_psrc_1 == io_writebackSignal_4),{(queue_3_psrc_1 == io_writebackSignal_3),{_zz_updatedEntry_3_srcReady_1,{_zz_updatedEntry_3_srcReady_1_1,_zz_updatedEntry_3_srcReady_1_2}}}})) || ((|{((queue_3_psrc_1 == io_earlyWakeup_7_payload) && io_earlyWakeup_7_valid),{(_zz_updatedEntry_3_srcReady_1_3 && io_earlyWakeup_6_valid),{_zz_updatedEntry_3_srcReady_1_4,{_zz_updatedEntry_3_srcReady_1_5,_zz_updatedEntry_3_srcReady_1_6}}}}) || ((queue_3_psrc_1 == io_wakeOut_payload) && io_wakeOut_valid)));
  end

  always @(*) begin
    shiftAhead[0] = ((|readyToIssue[0 : 0]) && io_output_ready);
    shiftAhead[1] = ((|readyToIssue[1 : 0]) && io_output_ready);
    shiftAhead[2] = ((|readyToIssue[2 : 0]) && io_output_ready);
    shiftAhead[3] = ((|readyToIssue[3 : 0]) && io_output_ready);
  end

  assign when_IssueQueue_l81 = shiftAhead[0];
  assign when_IssueQueue_l83 = writeVector[1];
  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_valid = appendEntry_valid;
      end else begin
        queueNext_0_valid = queue_1_valid;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_valid = appendEntry_valid;
      end else begin
        queueNext_0_valid = queue_0_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_0_robIdx = queue_1_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_0_robIdx = queue_0_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_0_branchInfo_predictPC = queue_1_branchInfo_predictPC;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_0_branchInfo_predictPC = queue_0_branchInfo_predictPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_0_branchInfo_predictResult = queue_1_branchInfo_predictResult;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_0_branchInfo_predictResult = queue_0_branchInfo_predictResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_0_exceptionInfo_exception = queue_1_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_0_exceptionInfo_exception = queue_0_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_0_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_0_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_0_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_0_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_pc = appendEntry_pc;
      end else begin
        queueNext_0_pc = queue_1_pc;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_pc = appendEntry_pc;
      end else begin
        queueNext_0_pc = queue_0_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_prd = appendEntry_prd;
      end else begin
        queueNext_0_prd = queue_1_prd;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_prd = appendEntry_prd;
      end else begin
        queueNext_0_prd = queue_0_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_0_psrc_0 = queue_1_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_0_psrc_0 = queue_0_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_0_psrc_1 = queue_1_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_0_psrc_1 = queue_0_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_imm = appendEntry_imm;
      end else begin
        queueNext_0_imm = queue_1_imm;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_imm = appendEntry_imm;
      end else begin
        queueNext_0_imm = queue_0_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_0_uop_aluOp = queue_1_uop_aluOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_0_uop_aluOp = queue_0_uop_aluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_0_uop_bruOp = queue_1_uop_bruOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_0_uop_bruOp = queue_0_uop_bruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_uop_cruOp = appendEntry_uop_cruOp;
      end else begin
        queueNext_0_uop_cruOp = queue_1_uop_cruOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_uop_cruOp = appendEntry_uop_cruOp;
      end else begin
        queueNext_0_uop_cruOp = queue_0_uop_cruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_0_roop_aluROOp = queue_1_roop_aluROOp;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_0_roop_aluROOp = queue_0_roop_aluROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_0_srcReady_0 = queue_1_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_0_srcReady_0 = queue_0_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81) begin
      if(when_IssueQueue_l83) begin
        queueNext_0_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_0_srcReady_1 = queue_1_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96) begin
        queueNext_0_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_0_srcReady_1 = queue_0_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96 = writeVector[0];
  assign when_IssueQueue_l81_1 = shiftAhead[1];
  assign when_IssueQueue_l83_1 = writeVector[2];
  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_valid = appendEntry_valid;
      end else begin
        queueNext_1_valid = queue_2_valid;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_valid = appendEntry_valid;
      end else begin
        queueNext_1_valid = queue_1_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_1_robIdx = queue_2_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_1_robIdx = queue_1_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_1_branchInfo_predictPC = queue_2_branchInfo_predictPC;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_1_branchInfo_predictPC = queue_1_branchInfo_predictPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_1_branchInfo_predictResult = queue_2_branchInfo_predictResult;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_1_branchInfo_predictResult = queue_1_branchInfo_predictResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_1_exceptionInfo_exception = queue_2_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_1_exceptionInfo_exception = queue_1_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_1_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_1_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_1_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_1_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_pc = appendEntry_pc;
      end else begin
        queueNext_1_pc = queue_2_pc;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_pc = appendEntry_pc;
      end else begin
        queueNext_1_pc = queue_1_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_prd = appendEntry_prd;
      end else begin
        queueNext_1_prd = queue_2_prd;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_prd = appendEntry_prd;
      end else begin
        queueNext_1_prd = queue_1_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_1_psrc_0 = queue_2_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_1_psrc_0 = queue_1_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_1_psrc_1 = queue_2_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_1_psrc_1 = queue_1_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_imm = appendEntry_imm;
      end else begin
        queueNext_1_imm = queue_2_imm;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_imm = appendEntry_imm;
      end else begin
        queueNext_1_imm = queue_1_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_1_uop_aluOp = queue_2_uop_aluOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_1_uop_aluOp = queue_1_uop_aluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_1_uop_bruOp = queue_2_uop_bruOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_1_uop_bruOp = queue_1_uop_bruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_uop_cruOp = appendEntry_uop_cruOp;
      end else begin
        queueNext_1_uop_cruOp = queue_2_uop_cruOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_uop_cruOp = appendEntry_uop_cruOp;
      end else begin
        queueNext_1_uop_cruOp = queue_1_uop_cruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_1_roop_aluROOp = queue_2_roop_aluROOp;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_1_roop_aluROOp = queue_1_roop_aluROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_1_srcReady_0 = queue_2_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_1_srcReady_0 = queue_1_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_1) begin
      if(when_IssueQueue_l83_1) begin
        queueNext_1_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_1_srcReady_1 = queue_2_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96_1) begin
        queueNext_1_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_1_srcReady_1 = queue_1_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_1 = writeVector[1];
  assign when_IssueQueue_l81_2 = shiftAhead[2];
  assign when_IssueQueue_l83_2 = writeVector[3];
  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_valid = appendEntry_valid;
      end else begin
        queueNext_2_valid = queue_3_valid;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_valid = appendEntry_valid;
      end else begin
        queueNext_2_valid = queue_2_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_2_robIdx = queue_3_robIdx;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_2_robIdx = queue_2_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_2_branchInfo_predictPC = queue_3_branchInfo_predictPC;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_2_branchInfo_predictPC = queue_2_branchInfo_predictPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_2_branchInfo_predictResult = queue_3_branchInfo_predictResult;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_2_branchInfo_predictResult = queue_2_branchInfo_predictResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_2_exceptionInfo_exception = queue_3_exceptionInfo_exception;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_2_exceptionInfo_exception = queue_2_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_2_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_2_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_2_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_2_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_pc = appendEntry_pc;
      end else begin
        queueNext_2_pc = queue_3_pc;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_pc = appendEntry_pc;
      end else begin
        queueNext_2_pc = queue_2_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_prd = appendEntry_prd;
      end else begin
        queueNext_2_prd = queue_3_prd;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_prd = appendEntry_prd;
      end else begin
        queueNext_2_prd = queue_2_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_2_psrc_0 = queue_3_psrc_0;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_2_psrc_0 = queue_2_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_2_psrc_1 = queue_3_psrc_1;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_2_psrc_1 = queue_2_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_imm = appendEntry_imm;
      end else begin
        queueNext_2_imm = queue_3_imm;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_imm = appendEntry_imm;
      end else begin
        queueNext_2_imm = queue_2_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_2_uop_aluOp = queue_3_uop_aluOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_2_uop_aluOp = queue_2_uop_aluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_2_uop_bruOp = queue_3_uop_bruOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_2_uop_bruOp = queue_2_uop_bruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_uop_cruOp = appendEntry_uop_cruOp;
      end else begin
        queueNext_2_uop_cruOp = queue_3_uop_cruOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_uop_cruOp = appendEntry_uop_cruOp;
      end else begin
        queueNext_2_uop_cruOp = queue_2_uop_cruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_2_roop_aluROOp = queue_3_roop_aluROOp;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_2_roop_aluROOp = queue_2_roop_aluROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_2_srcReady_0 = queue_3_srcReady_0;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_2_srcReady_0 = queue_2_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_2) begin
      if(when_IssueQueue_l83_2) begin
        queueNext_2_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_2_srcReady_1 = queue_3_srcReady_1;
      end
    end else begin
      if(when_IssueQueue_l96_2) begin
        queueNext_2_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_2_srcReady_1 = queue_2_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_2 = writeVector[2];
  assign when_IssueQueue_l81_3 = shiftAhead[3];
  assign when_IssueQueue_l89 = writeVector[4];
  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_valid = appendEntry_valid;
      end else begin
        queueNext_3_valid = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_valid = appendEntry_valid;
      end else begin
        queueNext_3_valid = queue_3_valid;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_3_robIdx = 5'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_robIdx = appendEntry_robIdx;
      end else begin
        queueNext_3_robIdx = queue_3_robIdx;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_3_branchInfo_predictPC = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchInfo_predictPC = appendEntry_branchInfo_predictPC;
      end else begin
        queueNext_3_branchInfo_predictPC = queue_3_branchInfo_predictPC;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_3_branchInfo_predictResult = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_branchInfo_predictResult = appendEntry_branchInfo_predictResult;
      end else begin
        queueNext_3_branchInfo_predictResult = queue_3_branchInfo_predictResult;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_3_exceptionInfo_exception = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_exception = appendEntry_exceptionInfo_exception;
      end else begin
        queueNext_3_exceptionInfo_exception = queue_3_exceptionInfo_exception;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_3_exceptionInfo_eCode = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_eCode = appendEntry_exceptionInfo_eCode;
      end else begin
        queueNext_3_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_3_exceptionInfo_eSubCode = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_exceptionInfo_eSubCode = appendEntry_exceptionInfo_eSubCode;
      end else begin
        queueNext_3_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_pc = appendEntry_pc;
      end else begin
        queueNext_3_pc = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_pc = appendEntry_pc;
      end else begin
        queueNext_3_pc = queue_3_pc;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_prd = appendEntry_prd;
      end else begin
        queueNext_3_prd = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_prd = appendEntry_prd;
      end else begin
        queueNext_3_prd = queue_3_prd;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_3_psrc_0 = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_psrc_0 = appendEntry_psrc_0;
      end else begin
        queueNext_3_psrc_0 = queue_3_psrc_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_3_psrc_1 = 6'h00;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_psrc_1 = appendEntry_psrc_1;
      end else begin
        queueNext_3_psrc_1 = queue_3_psrc_1;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_imm = appendEntry_imm;
      end else begin
        queueNext_3_imm = 32'h00000000;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_imm = appendEntry_imm;
      end else begin
        queueNext_3_imm = queue_3_imm;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_3_uop_aluOp = ALUOp_add;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_uop_aluOp = appendEntry_uop_aluOp;
      end else begin
        queueNext_3_uop_aluOp = queue_3_uop_aluOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_3_uop_bruOp = BRUOp_nop;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_uop_bruOp = appendEntry_uop_bruOp;
      end else begin
        queueNext_3_uop_bruOp = queue_3_uop_bruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_uop_cruOp = appendEntry_uop_cruOp;
      end else begin
        queueNext_3_uop_cruOp = CRUOp_nop;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_uop_cruOp = appendEntry_uop_cruOp;
      end else begin
        queueNext_3_uop_cruOp = queue_3_uop_cruOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_3_roop_aluROOp = ALUROOp_reg_1;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_roop_aluROOp = appendEntry_roop_aluROOp;
      end else begin
        queueNext_3_roop_aluROOp = queue_3_roop_aluROOp;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_3_srcReady_0 = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_srcReady_0 = appendEntry_srcReady_0;
      end else begin
        queueNext_3_srcReady_0 = queue_3_srcReady_0;
      end
    end
  end

  always @(*) begin
    if(when_IssueQueue_l81_3) begin
      if(when_IssueQueue_l89) begin
        queueNext_3_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_3_srcReady_1 = 1'b0;
      end
    end else begin
      if(when_IssueQueue_l96_3) begin
        queueNext_3_srcReady_1 = appendEntry_srcReady_1;
      end else begin
        queueNext_3_srcReady_1 = queue_3_srcReady_1;
      end
    end
  end

  assign when_IssueQueue_l96_3 = writeVector[3];
  always @(*) begin
    _zz_io_csrInQueue[0] = ((queue_0_roop_aluROOp == ALUROOp_csr) && queue_0_valid);
    _zz_io_csrInQueue[1] = ((queue_1_roop_aluROOp == ALUROOp_csr) && queue_1_valid);
    _zz_io_csrInQueue[2] = ((queue_2_roop_aluROOp == ALUROOp_csr) && queue_2_valid);
    _zz_io_csrInQueue[3] = ((queue_3_roop_aluROOp == ALUROOp_csr) && queue_3_valid);
  end

  assign io_csrInQueue = (|_zz_io_csrInQueue);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_input_ready = ((|emptyEntry[3 : 0]) || io_output_fire);
  assign _zz_issueEntry_valid = issueVector[3];
  assign _zz_issueEntry_valid_1 = (issueVector[1] || _zz_issueEntry_valid);
  assign _zz_issueEntry_valid_2 = (issueVector[2] || _zz_issueEntry_valid);
  assign _zz_issueEntry_valid_3 = {_zz_issueEntry_valid_2,_zz_issueEntry_valid_1};
  assign issueEntry_valid = _zz_issueEntry_valid_4;
  assign issueEntry_robIdx = _zz_issueEntry_robIdx;
  assign issueEntry_branchInfo_predictPC = _zz_issueEntry_branchInfo_predictPC;
  assign issueEntry_branchInfo_predictResult = _zz_issueEntry_branchInfo_predictResult;
  assign issueEntry_exceptionInfo_exception = _zz_issueEntry_exceptionInfo_exception;
  assign issueEntry_exceptionInfo_eCode = _zz_issueEntry_exceptionInfo_eCode;
  assign issueEntry_exceptionInfo_eSubCode = _zz_issueEntry_exceptionInfo_eSubCode;
  assign issueEntry_pc = _zz_issueEntry_pc;
  assign issueEntry_prd = _zz_issueEntry_prd;
  assign issueEntry_psrc_0 = _zz_issueEntry_psrc_0;
  assign issueEntry_psrc_1 = _zz_issueEntry_psrc_1;
  assign issueEntry_imm = _zz_issueEntry_imm;
  assign issueEntry_uop_aluOp = _zz_issueEntry_uop_aluOp;
  assign issueEntry_uop_bruOp = _zz_issueEntry_uop_bruOp;
  assign issueEntry_uop_cruOp = _zz_issueEntry_uop_cruOp;
  assign issueEntry_roop_aluROOp = _zz_issueEntry_roop_aluROOp;
  assign issueEntry_srcReady_0 = _zz_issueEntry_srcReady_0;
  assign issueEntry_srcReady_1 = _zz_issueEntry_srcReady_1;
  assign io_output_valid = (|readyToIssue);
  assign io_output_payload_robIdx = issueEntry_robIdx;
  assign io_output_payload_branchInfo_predictPC = issueEntry_branchInfo_predictPC;
  assign io_output_payload_branchInfo_predictResult = issueEntry_branchInfo_predictResult;
  assign io_output_payload_exceptionInfo_exception = issueEntry_exceptionInfo_exception;
  assign io_output_payload_exceptionInfo_eCode = issueEntry_exceptionInfo_eCode;
  assign io_output_payload_exceptionInfo_eSubCode = issueEntry_exceptionInfo_eSubCode;
  assign io_output_payload_pc = issueEntry_pc;
  assign io_output_payload_prd = issueEntry_prd;
  assign io_output_payload_psrc_0 = issueEntry_psrc_0;
  assign io_output_payload_psrc_1 = issueEntry_psrc_1;
  assign io_output_payload_imm = issueEntry_imm;
  assign io_output_payload_uop_aluOp = issueEntry_uop_aluOp;
  assign io_output_payload_uop_bruOp = issueEntry_uop_bruOp;
  assign io_output_payload_uop_cruOp = issueEntry_uop_cruOp;
  assign io_output_payload_roop_aluROOp = issueEntry_roop_aluROOp;
  assign io_wakeOut_payload = issueEntry_prd;
  assign io_wakeOut_valid = io_output_fire;
  always @(posedge aclk) begin
    if(!cpuClockingArea_areaFlushReset_newReset) begin
      queue_0_valid <= 1'b0;
      queue_0_robIdx <= 5'h00;
      queue_0_branchInfo_predictPC <= 32'h00000000;
      queue_0_branchInfo_predictResult <= 1'b0;
      queue_0_exceptionInfo_exception <= 1'b0;
      queue_0_exceptionInfo_eCode <= 6'h00;
      queue_0_exceptionInfo_eSubCode <= 1'b0;
      queue_0_pc <= 32'h00000000;
      queue_0_prd <= 6'h00;
      queue_0_psrc_0 <= 6'h00;
      queue_0_psrc_1 <= 6'h00;
      queue_0_imm <= 32'h00000000;
      queue_0_uop_aluOp <= ALUOp_add;
      queue_0_uop_bruOp <= BRUOp_nop;
      queue_0_uop_cruOp <= CRUOp_nop;
      queue_0_roop_aluROOp <= ALUROOp_reg_1;
      queue_0_srcReady_0 <= 1'b0;
      queue_0_srcReady_1 <= 1'b0;
      queue_1_valid <= 1'b0;
      queue_1_robIdx <= 5'h00;
      queue_1_branchInfo_predictPC <= 32'h00000000;
      queue_1_branchInfo_predictResult <= 1'b0;
      queue_1_exceptionInfo_exception <= 1'b0;
      queue_1_exceptionInfo_eCode <= 6'h00;
      queue_1_exceptionInfo_eSubCode <= 1'b0;
      queue_1_pc <= 32'h00000000;
      queue_1_prd <= 6'h00;
      queue_1_psrc_0 <= 6'h00;
      queue_1_psrc_1 <= 6'h00;
      queue_1_imm <= 32'h00000000;
      queue_1_uop_aluOp <= ALUOp_add;
      queue_1_uop_bruOp <= BRUOp_nop;
      queue_1_uop_cruOp <= CRUOp_nop;
      queue_1_roop_aluROOp <= ALUROOp_reg_1;
      queue_1_srcReady_0 <= 1'b0;
      queue_1_srcReady_1 <= 1'b0;
      queue_2_valid <= 1'b0;
      queue_2_robIdx <= 5'h00;
      queue_2_branchInfo_predictPC <= 32'h00000000;
      queue_2_branchInfo_predictResult <= 1'b0;
      queue_2_exceptionInfo_exception <= 1'b0;
      queue_2_exceptionInfo_eCode <= 6'h00;
      queue_2_exceptionInfo_eSubCode <= 1'b0;
      queue_2_pc <= 32'h00000000;
      queue_2_prd <= 6'h00;
      queue_2_psrc_0 <= 6'h00;
      queue_2_psrc_1 <= 6'h00;
      queue_2_imm <= 32'h00000000;
      queue_2_uop_aluOp <= ALUOp_add;
      queue_2_uop_bruOp <= BRUOp_nop;
      queue_2_uop_cruOp <= CRUOp_nop;
      queue_2_roop_aluROOp <= ALUROOp_reg_1;
      queue_2_srcReady_0 <= 1'b0;
      queue_2_srcReady_1 <= 1'b0;
      queue_3_valid <= 1'b0;
      queue_3_robIdx <= 5'h00;
      queue_3_branchInfo_predictPC <= 32'h00000000;
      queue_3_branchInfo_predictResult <= 1'b0;
      queue_3_exceptionInfo_exception <= 1'b0;
      queue_3_exceptionInfo_eCode <= 6'h00;
      queue_3_exceptionInfo_eSubCode <= 1'b0;
      queue_3_pc <= 32'h00000000;
      queue_3_prd <= 6'h00;
      queue_3_psrc_0 <= 6'h00;
      queue_3_psrc_1 <= 6'h00;
      queue_3_imm <= 32'h00000000;
      queue_3_uop_aluOp <= ALUOp_add;
      queue_3_uop_bruOp <= BRUOp_nop;
      queue_3_uop_cruOp <= CRUOp_nop;
      queue_3_roop_aluROOp <= ALUROOp_reg_1;
      queue_3_srcReady_0 <= 1'b0;
      queue_3_srcReady_1 <= 1'b0;
    end else begin
      queue_0_valid <= queueNext_0_valid;
      queue_0_robIdx <= queueNext_0_robIdx;
      queue_0_branchInfo_predictPC <= queueNext_0_branchInfo_predictPC;
      queue_0_branchInfo_predictResult <= queueNext_0_branchInfo_predictResult;
      queue_0_exceptionInfo_exception <= queueNext_0_exceptionInfo_exception;
      queue_0_exceptionInfo_eCode <= queueNext_0_exceptionInfo_eCode;
      queue_0_exceptionInfo_eSubCode <= queueNext_0_exceptionInfo_eSubCode;
      queue_0_pc <= queueNext_0_pc;
      queue_0_prd <= queueNext_0_prd;
      queue_0_psrc_0 <= queueNext_0_psrc_0;
      queue_0_psrc_1 <= queueNext_0_psrc_1;
      queue_0_imm <= queueNext_0_imm;
      queue_0_uop_aluOp <= queueNext_0_uop_aluOp;
      queue_0_uop_bruOp <= queueNext_0_uop_bruOp;
      queue_0_uop_cruOp <= queueNext_0_uop_cruOp;
      queue_0_roop_aluROOp <= queueNext_0_roop_aluROOp;
      queue_0_srcReady_0 <= queueNext_0_srcReady_0;
      queue_0_srcReady_1 <= queueNext_0_srcReady_1;
      queue_1_valid <= queueNext_1_valid;
      queue_1_robIdx <= queueNext_1_robIdx;
      queue_1_branchInfo_predictPC <= queueNext_1_branchInfo_predictPC;
      queue_1_branchInfo_predictResult <= queueNext_1_branchInfo_predictResult;
      queue_1_exceptionInfo_exception <= queueNext_1_exceptionInfo_exception;
      queue_1_exceptionInfo_eCode <= queueNext_1_exceptionInfo_eCode;
      queue_1_exceptionInfo_eSubCode <= queueNext_1_exceptionInfo_eSubCode;
      queue_1_pc <= queueNext_1_pc;
      queue_1_prd <= queueNext_1_prd;
      queue_1_psrc_0 <= queueNext_1_psrc_0;
      queue_1_psrc_1 <= queueNext_1_psrc_1;
      queue_1_imm <= queueNext_1_imm;
      queue_1_uop_aluOp <= queueNext_1_uop_aluOp;
      queue_1_uop_bruOp <= queueNext_1_uop_bruOp;
      queue_1_uop_cruOp <= queueNext_1_uop_cruOp;
      queue_1_roop_aluROOp <= queueNext_1_roop_aluROOp;
      queue_1_srcReady_0 <= queueNext_1_srcReady_0;
      queue_1_srcReady_1 <= queueNext_1_srcReady_1;
      queue_2_valid <= queueNext_2_valid;
      queue_2_robIdx <= queueNext_2_robIdx;
      queue_2_branchInfo_predictPC <= queueNext_2_branchInfo_predictPC;
      queue_2_branchInfo_predictResult <= queueNext_2_branchInfo_predictResult;
      queue_2_exceptionInfo_exception <= queueNext_2_exceptionInfo_exception;
      queue_2_exceptionInfo_eCode <= queueNext_2_exceptionInfo_eCode;
      queue_2_exceptionInfo_eSubCode <= queueNext_2_exceptionInfo_eSubCode;
      queue_2_pc <= queueNext_2_pc;
      queue_2_prd <= queueNext_2_prd;
      queue_2_psrc_0 <= queueNext_2_psrc_0;
      queue_2_psrc_1 <= queueNext_2_psrc_1;
      queue_2_imm <= queueNext_2_imm;
      queue_2_uop_aluOp <= queueNext_2_uop_aluOp;
      queue_2_uop_bruOp <= queueNext_2_uop_bruOp;
      queue_2_uop_cruOp <= queueNext_2_uop_cruOp;
      queue_2_roop_aluROOp <= queueNext_2_roop_aluROOp;
      queue_2_srcReady_0 <= queueNext_2_srcReady_0;
      queue_2_srcReady_1 <= queueNext_2_srcReady_1;
      queue_3_valid <= queueNext_3_valid;
      queue_3_robIdx <= queueNext_3_robIdx;
      queue_3_branchInfo_predictPC <= queueNext_3_branchInfo_predictPC;
      queue_3_branchInfo_predictResult <= queueNext_3_branchInfo_predictResult;
      queue_3_exceptionInfo_exception <= queueNext_3_exceptionInfo_exception;
      queue_3_exceptionInfo_eCode <= queueNext_3_exceptionInfo_eCode;
      queue_3_exceptionInfo_eSubCode <= queueNext_3_exceptionInfo_eSubCode;
      queue_3_pc <= queueNext_3_pc;
      queue_3_prd <= queueNext_3_prd;
      queue_3_psrc_0 <= queueNext_3_psrc_0;
      queue_3_psrc_1 <= queueNext_3_psrc_1;
      queue_3_imm <= queueNext_3_imm;
      queue_3_uop_aluOp <= queueNext_3_uop_aluOp;
      queue_3_uop_bruOp <= queueNext_3_uop_bruOp;
      queue_3_uop_cruOp <= queueNext_3_uop_cruOp;
      queue_3_roop_aluROOp <= queueNext_3_roop_aluROOp;
      queue_3_srcReady_0 <= queueNext_3_srcReady_0;
      queue_3_srcReady_1 <= queueNext_3_srcReady_1;
    end
  end


endmodule

module Dispatcher (
  output wire [1:0]    io_input_allowMask,
  input  wire [1:0]    io_input_availMask,
  input  wire [31:0]   io_input_info_0_inst,
  input  wire [31:0]   io_input_info_0_branchInfo_predictPC,
  input  wire          io_input_info_0_branchInfo_predictResult,
  input  wire          io_input_info_0_exceptionInfo_exception,
  input  wire [5:0]    io_input_info_0_exceptionInfo_eCode,
  input  wire [0:0]    io_input_info_0_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_info_0_pc,
  input  wire [31:0]   io_input_info_1_inst,
  input  wire [31:0]   io_input_info_1_branchInfo_predictPC,
  input  wire          io_input_info_1_branchInfo_predictResult,
  input  wire          io_input_info_1_exceptionInfo_exception,
  input  wire [5:0]    io_input_info_1_exceptionInfo_eCode,
  input  wire [0:0]    io_input_info_1_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_info_1_pc,
  input  wire [2:0]    io_input_dispatchInfo_0_fuType,
  input  wire [4:0]    io_input_dispatchInfo_0_ard,
  input  wire [4:0]    io_input_dispatchInfo_0_asrc_0,
  input  wire [4:0]    io_input_dispatchInfo_0_asrc_1,
  input  wire [2:0]    io_input_dispatchInfo_1_fuType,
  input  wire [4:0]    io_input_dispatchInfo_1_ard,
  input  wire [4:0]    io_input_dispatchInfo_1_asrc_0,
  input  wire [4:0]    io_input_dispatchInfo_1_asrc_1,
  input  wire          io_aluHasCSRInst_0,
  input  wire          io_aluHasCSRInst_1,
  output wire [1:0]    io_rob_allowMask,
  input  wire [1:0]    io_rob_availMask,
  input  wire [4:0]    io_rob_robIdx_0,
  input  wire [4:0]    io_rob_robIdx_1,
  output wire [31:0]   io_rob_pc_0,
  output wire [31:0]   io_rob_pc_1,
  output wire [4:0]    io_rob_ard_0,
  output wire [4:0]    io_rob_ard_1,
  output wire [5:0]    io_rob_prd_0,
  output wire [5:0]    io_rob_prd_1,
  output wire [5:0]    io_rob_pprd_0,
  output wire [5:0]    io_rob_pprd_1,
  output wire [3:0]    io_rob_specialOp_0,
  output wire [3:0]    io_rob_specialOp_1,
  output wire [4:0]    io_sratWrite_0_ard,
  output wire [5:0]    io_sratWrite_0_prd,
  output wire          io_sratWrite_0_wen,
  output wire [4:0]    io_sratWrite_1_ard,
  output wire [5:0]    io_sratWrite_1_prd,
  output wire          io_sratWrite_1_wen,
  output wire [4:0]    io_sratReadSrc_0_0_ard,
  input  wire [5:0]    io_sratReadSrc_0_0_prd,
  input  wire          io_sratReadSrc_0_0_valid,
  output wire [4:0]    io_sratReadSrc_0_1_ard,
  input  wire [5:0]    io_sratReadSrc_0_1_prd,
  input  wire          io_sratReadSrc_0_1_valid,
  output wire [4:0]    io_sratReadSrc_1_0_ard,
  input  wire [5:0]    io_sratReadSrc_1_0_prd,
  input  wire          io_sratReadSrc_1_0_valid,
  output wire [4:0]    io_sratReadSrc_1_1_ard,
  input  wire [5:0]    io_sratReadSrc_1_1_prd,
  input  wire          io_sratReadSrc_1_1_valid,
  output wire [4:0]    io_sratReadPPRD_0_ard,
  input  wire [5:0]    io_sratReadPPRD_0_prd,
  input  wire          io_sratReadPPRD_0_valid,
  output wire [4:0]    io_sratReadPPRD_1_ard,
  input  wire [5:0]    io_sratReadPPRD_1_prd,
  input  wire          io_sratReadPPRD_1_valid,
  output wire [1:0]    io_freelist_disPatchNum,
  input  wire [1:0]    io_freelist_availMask,
  input  wire [5:0]    io_freelist_prfIdx_0,
  input  wire [5:0]    io_freelist_prfIdx_1,
  input  wire [1:0]    _zz_when_Decoder_l40,
  output wire          io_alu0IQ_valid,
  input  wire          io_alu0IQ_ready,
  output wire [4:0]    io_alu0IQ_payload_robIdx,
  output wire [31:0]   io_alu0IQ_payload_branchInfo_predictPC,
  output wire          io_alu0IQ_payload_branchInfo_predictResult,
  output wire          io_alu0IQ_payload_exceptionInfo_exception,
  output wire [5:0]    io_alu0IQ_payload_exceptionInfo_eCode,
  output wire [0:0]    io_alu0IQ_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_alu0IQ_payload_pc,
  output wire [5:0]    io_alu0IQ_payload_prd,
  output wire [5:0]    io_alu0IQ_payload_psrc_0,
  output wire [5:0]    io_alu0IQ_payload_psrc_1,
  output wire [31:0]   io_alu0IQ_payload_imm,
  output wire [3:0]    io_alu0IQ_payload_uop_aluOp,
  output wire [1:0]    io_alu0IQ_payload_uop_bruOp,
  output wire [1:0]    io_alu0IQ_payload_uop_cruOp,
  output wire [2:0]    io_alu0IQ_payload_roop_aluROOp,
  output wire          io_alu0IQ_payload_srcReady_0,
  output wire          io_alu0IQ_payload_srcReady_1,
  output wire          io_alu1IQ_valid,
  input  wire          io_alu1IQ_ready,
  output wire [4:0]    io_alu1IQ_payload_robIdx,
  output wire [31:0]   io_alu1IQ_payload_branchInfo_predictPC,
  output wire          io_alu1IQ_payload_branchInfo_predictResult,
  output wire          io_alu1IQ_payload_exceptionInfo_exception,
  output wire [5:0]    io_alu1IQ_payload_exceptionInfo_eCode,
  output wire [0:0]    io_alu1IQ_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_alu1IQ_payload_pc,
  output wire [5:0]    io_alu1IQ_payload_prd,
  output wire [5:0]    io_alu1IQ_payload_psrc_0,
  output wire [5:0]    io_alu1IQ_payload_psrc_1,
  output wire [31:0]   io_alu1IQ_payload_imm,
  output wire [3:0]    io_alu1IQ_payload_uop_aluOp,
  output wire [1:0]    io_alu1IQ_payload_uop_bruOp,
  output wire [2:0]    io_alu1IQ_payload_roop_aluROOp,
  output wire [1:0]    io_alu1IQ_payload_roop_cruROOp,
  output wire          io_alu1IQ_payload_srcReady_0,
  output wire          io_alu1IQ_payload_srcReady_1,
  output wire          io_muluIQ_valid,
  input  wire          io_muluIQ_ready,
  output wire [4:0]    io_muluIQ_payload_robIdx,
  output wire [31:0]   io_muluIQ_payload_branchResult_targetPC,
  output wire          io_muluIQ_payload_branchResult_branchResult,
  output wire          io_muluIQ_payload_branchResult_predictFail,
  output wire          io_muluIQ_payload_exceptionInfo_exception,
  output wire [5:0]    io_muluIQ_payload_exceptionInfo_eCode,
  output wire [0:0]    io_muluIQ_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_muluIQ_payload_pc,
  output wire [5:0]    io_muluIQ_payload_prd,
  output wire [5:0]    io_muluIQ_payload_psrc_0,
  output wire [5:0]    io_muluIQ_payload_psrc_1,
  output wire [31:0]   io_muluIQ_payload_imm,
  output wire [1:0]    io_muluIQ_payload_uop_muluOp,
  output wire          io_muluIQ_payload_srcReady_0,
  output wire          io_muluIQ_payload_srcReady_1,
  output wire          io_divuIQ_valid,
  input  wire          io_divuIQ_ready,
  output wire [4:0]    io_divuIQ_payload_robIdx,
  output wire [31:0]   io_divuIQ_payload_branchResult_targetPC,
  output wire          io_divuIQ_payload_branchResult_branchResult,
  output wire          io_divuIQ_payload_branchResult_predictFail,
  output wire          io_divuIQ_payload_exceptionInfo_exception,
  output wire [5:0]    io_divuIQ_payload_exceptionInfo_eCode,
  output wire [0:0]    io_divuIQ_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_divuIQ_payload_pc,
  output wire [5:0]    io_divuIQ_payload_prd,
  output wire [5:0]    io_divuIQ_payload_psrc_0,
  output wire [5:0]    io_divuIQ_payload_psrc_1,
  output wire [31:0]   io_divuIQ_payload_imm,
  output wire [1:0]    io_divuIQ_payload_uop_divuOp,
  output wire          io_divuIQ_payload_srcReady_0,
  output wire          io_divuIQ_payload_srcReady_1,
  output wire          io_lsuIQ_valid,
  input  wire          io_lsuIQ_ready,
  output wire [4:0]    io_lsuIQ_payload_robIdx,
  output wire [31:0]   io_lsuIQ_payload_branchResult_targetPC,
  output wire          io_lsuIQ_payload_branchResult_branchResult,
  output wire          io_lsuIQ_payload_branchResult_predictFail,
  output wire          io_lsuIQ_payload_exceptionInfo_exception,
  output wire [5:0]    io_lsuIQ_payload_exceptionInfo_eCode,
  output wire [0:0]    io_lsuIQ_payload_exceptionInfo_eSubCode,
  output wire [31:0]   io_lsuIQ_payload_pc,
  output wire [5:0]    io_lsuIQ_payload_prd,
  output wire [5:0]    io_lsuIQ_payload_psrc_0,
  output wire [5:0]    io_lsuIQ_payload_psrc_1,
  output wire [31:0]   io_lsuIQ_payload_imm,
  output wire [3:0]    io_lsuIQ_payload_uop_lsuOp,
  output wire [4:0]    io_lsuIQ_payload_uop_lsuCoOp,
  output wire [0:0]    io_lsuIQ_payload_roop_lsuROOp,
  output wire          io_lsuIQ_payload_srcReady_0,
  output wire          io_lsuIQ_payload_srcReady_1
);
  localparam FUType_alu = 3'd0;
  localparam FUType_csr = 3'd1;
  localparam FUType_counter = 3'd2;
  localparam FUType_lsu = 3'd3;
  localparam FUType_mulu = 3'd4;
  localparam FUType_divu = 3'd5;
  localparam ROBSpecialOp_nop = 4'd0;
  localparam ROBSpecialOp_bpuUpdate = 4'd1;
  localparam ROBSpecialOp_lsuAction = 4'd2;
  localparam ROBSpecialOp_ll = 4'd3;
  localparam ROBSpecialOp_writeCSR = 4'd4;
  localparam ROBSpecialOp_ertn = 4'd5;
  localparam ROBSpecialOp_idle = 4'd6;
  localparam ROBSpecialOp_readCSR = 4'd7;
  localparam ROBSpecialOp_readCNT = 4'd8;
  localparam ALUOp_add = 4'd0;
  localparam ALUOp_sub = 4'd1;
  localparam ALUOp_slt = 4'd2;
  localparam ALUOp_sltu = 4'd3;
  localparam ALUOp_eq = 4'd4;
  localparam ALUOp_nor_1 = 4'd5;
  localparam ALUOp_and_1 = 4'd6;
  localparam ALUOp_or_1 = 4'd7;
  localparam ALUOp_xor_1 = 4'd8;
  localparam ALUOp_sll_1 = 4'd9;
  localparam ALUOp_srl_1 = 4'd10;
  localparam ALUOp_sra_1 = 4'd11;
  localparam ALUOp_passa = 4'd12;
  localparam ALUOp_passb = 4'd13;
  localparam BRUOp_nop = 2'd0;
  localparam BRUOp_add = 2'd1;
  localparam BRUOp_cadd = 2'd2;
  localparam BRUOp_ncadd = 2'd3;
  localparam CRUOp_nop = 2'd0;
  localparam CRUOp_pass = 2'd1;
  localparam CRUOp_mask = 2'd2;
  localparam ALUROOp_reg_1 = 3'd0;
  localparam ALUROOp_regimm = 3'd1;
  localparam ALUROOp_pcimm = 3'd2;
  localparam ALUROOp_csr = 3'd3;
  localparam ALUROOp_linkpc = 3'd4;
  localparam ALUROOp_linkreg = 3'd5;
  localparam CRUROOp_id = 2'd0;
  localparam CRUROOp_lo = 2'd1;
  localparam CRUROOp_hi = 2'd2;
  localparam MULUOp_mullo = 2'd0;
  localparam MULUOp_mulhi = 2'd1;
  localparam MULUOp_mulhiu = 2'd2;
  localparam DIVUOp_div = 2'd0;
  localparam DIVUOp_divu = 2'd1;
  localparam DIVUOp_mod_1 = 2'd2;
  localparam DIVUOp_modu = 2'd3;
  localparam LSUOp_cacop = 4'd0;
  localparam LSUOp_tlbsrch = 4'd1;
  localparam LSUOp_tlbrd = 4'd2;
  localparam LSUOp_tlbwr = 4'd3;
  localparam LSUOp_tlbfill = 4'd4;
  localparam LSUOp_invtlb = 4'd5;
  localparam LSUOp_ll = 4'd6;
  localparam LSUOp_sc = 4'd7;
  localparam LSUOp_ld = 4'd8;
  localparam LSUOp_ldu = 4'd9;
  localparam LSUOp_st = 4'd10;
  localparam LSUOp_preld = 4'd11;
  localparam LSUOp_dbar = 4'd12;
  localparam LSUOp_ibar = 4'd13;
  localparam LSUROOp_reg_1 = 1'd0;
  localparam LSUROOp_regimm = 1'd1;

  wire       [31:0]   decoder_0_io_branchInfo_predictPC;
  wire                decoder_0_io_branchInfo_predictResult;
  wire       [31:0]   decoder_0_io_branchResult_targetPC;
  wire                decoder_0_io_branchResult_branchResult;
  wire                decoder_0_io_branchResult_predictFail;
  wire                decoder_0_io_exceptionInfo_exception;
  wire       [5:0]    decoder_0_io_exceptionInfo_eCode;
  wire       [0:0]    decoder_0_io_exceptionInfo_eSubCode;
  wire       [31:0]   decoder_0_io_pc;
  wire       [3:0]    decoder_0_io_specialOp;
  wire       [31:0]   decoder_0_io_imm;
  wire       [3:0]    decoder_0_io_uopALU0_aluOp;
  wire       [1:0]    decoder_0_io_uopALU0_bruOp;
  wire       [1:0]    decoder_0_io_uopALU0_cruOp;
  wire       [3:0]    decoder_0_io_uopALU1_aluOp;
  wire       [1:0]    decoder_0_io_uopALU1_bruOp;
  wire       [1:0]    decoder_0_io_uopMULU_muluOp;
  wire       [1:0]    decoder_0_io_uopDIVU_divuOp;
  wire       [3:0]    decoder_0_io_uopLSU_lsuOp;
  wire       [4:0]    decoder_0_io_uopLSU_lsuCoOp;
  wire       [2:0]    decoder_0_io_roopALU0_aluROOp;
  wire       [2:0]    decoder_0_io_roopALU1_aluROOp;
  wire       [1:0]    decoder_0_io_roopALU1_cruROOp;
  wire       [0:0]    decoder_0_io_roopLSU_lsuROOp;
  wire       [31:0]   decoder_1_1_io_branchInfo_predictPC;
  wire                decoder_1_1_io_branchInfo_predictResult;
  wire       [31:0]   decoder_1_1_io_branchResult_targetPC;
  wire                decoder_1_1_io_branchResult_branchResult;
  wire                decoder_1_1_io_branchResult_predictFail;
  wire                decoder_1_1_io_exceptionInfo_exception;
  wire       [5:0]    decoder_1_1_io_exceptionInfo_eCode;
  wire       [0:0]    decoder_1_1_io_exceptionInfo_eSubCode;
  wire       [31:0]   decoder_1_1_io_pc;
  wire       [3:0]    decoder_1_1_io_specialOp;
  wire       [31:0]   decoder_1_1_io_imm;
  wire       [3:0]    decoder_1_1_io_uopALU0_aluOp;
  wire       [1:0]    decoder_1_1_io_uopALU0_bruOp;
  wire       [1:0]    decoder_1_1_io_uopALU0_cruOp;
  wire       [3:0]    decoder_1_1_io_uopALU1_aluOp;
  wire       [1:0]    decoder_1_1_io_uopALU1_bruOp;
  wire       [1:0]    decoder_1_1_io_uopMULU_muluOp;
  wire       [1:0]    decoder_1_1_io_uopDIVU_divuOp;
  wire       [3:0]    decoder_1_1_io_uopLSU_lsuOp;
  wire       [4:0]    decoder_1_1_io_uopLSU_lsuCoOp;
  wire       [2:0]    decoder_1_1_io_roopALU0_aluROOp;
  wire       [2:0]    decoder_1_1_io_roopALU1_aluROOp;
  wire       [1:0]    decoder_1_1_io_roopALU1_cruROOp;
  wire       [0:0]    decoder_1_1_io_roopLSU_lsuROOp;
  reg        [5:0]    _zz_freelistRdShuffle_1;
  reg        [0:0]    _zz_freelistRdShuffle_1_1;
  wire       [0:0]    _zz_freelistRdShuffle_1_2;
  reg        [0:0]    _zz_freelistAvail;
  wire       [0:0]    _zz_freelistAvail_1;
  wire       [1:0]    _zz_alu0Sel_1;
  wire       [1:0]    _zz_alu1Sel_1;
  wire       [1:0]    _zz_muluReq_ohFirst_masked;
  wire       [1:0]    _zz_divuReq_ohFirst_masked;
  wire       [1:0]    _zz_lsuReq_ohFirst_masked;
  reg        [1:0]    _zz_io_freelist_disPatchNum;
  wire       [1:0]    _zz_io_freelist_disPatchNum_1;
  wire       [1:0]    _zz__zz_actualSrc_1_0_2;
  wire       [1:0]    _zz__zz_actualSrc_1_1_2;
  wire       [1:0]    _zz__zz_actualpRd_1_3;
  wire       [1:0]    resAvail;
  reg        [1:0]    needRd;
  reg        [5:0]    freelistRdShuffle_0;
  reg        [5:0]    freelistRdShuffle_1;
  reg        [1:0]    freelistAvail;
  wire                when_Dispatcher_l34;
  wire                when_Dispatcher_l42;
  wire       [1:0]    iqAvail;
  reg        [1:0]    csrReq;
  reg        [1:0]    counterReq;
  reg        [1:0]    alu0Req;
  reg        [1:0]    alu1Req;
  reg        [1:0]    muluReq;
  reg        [1:0]    divuReq;
  reg        [1:0]    lsuReq;
  wire       [1:0]    _zz_alu0Sel;
  wire       [1:0]    alu0Sel;
  wire       [1:0]    _zz_alu1Sel;
  wire       [1:0]    alu1Sel;
  wire       [1:0]    muluReq_ohFirst_input;
  wire       [1:0]    muluReq_ohFirst_masked;
  wire       [1:0]    muluSel;
  wire       [1:0]    divuReq_ohFirst_input;
  wire       [1:0]    divuReq_ohFirst_masked;
  wire       [1:0]    divuSel;
  wire       [1:0]    lsuReq_ohFirst_input;
  wire       [1:0]    lsuReq_ohFirst_masked;
  wire       [1:0]    lsuSel;
  reg        [1:0]    dispatchMask;
  wire       [4:0]    alu0Candidate_0_robIdx;
  wire       [31:0]   alu0Candidate_0_branchInfo_predictPC;
  wire                alu0Candidate_0_branchInfo_predictResult;
  wire                alu0Candidate_0_exceptionInfo_exception;
  wire       [5:0]    alu0Candidate_0_exceptionInfo_eCode;
  wire       [0:0]    alu0Candidate_0_exceptionInfo_eSubCode;
  wire       [31:0]   alu0Candidate_0_pc;
  wire       [5:0]    alu0Candidate_0_prd;
  wire       [5:0]    alu0Candidate_0_psrc_0;
  wire       [5:0]    alu0Candidate_0_psrc_1;
  wire       [31:0]   alu0Candidate_0_imm;
  wire       [3:0]    alu0Candidate_0_uop_aluOp;
  wire       [1:0]    alu0Candidate_0_uop_bruOp;
  wire       [1:0]    alu0Candidate_0_uop_cruOp;
  wire       [2:0]    alu0Candidate_0_roop_aluROOp;
  wire                alu0Candidate_0_srcReady_0;
  wire                alu0Candidate_0_srcReady_1;
  wire       [4:0]    alu0Candidate_1_robIdx;
  wire       [31:0]   alu0Candidate_1_branchInfo_predictPC;
  wire                alu0Candidate_1_branchInfo_predictResult;
  wire                alu0Candidate_1_exceptionInfo_exception;
  wire       [5:0]    alu0Candidate_1_exceptionInfo_eCode;
  wire       [0:0]    alu0Candidate_1_exceptionInfo_eSubCode;
  wire       [31:0]   alu0Candidate_1_pc;
  wire       [5:0]    alu0Candidate_1_prd;
  wire       [5:0]    alu0Candidate_1_psrc_0;
  wire       [5:0]    alu0Candidate_1_psrc_1;
  wire       [31:0]   alu0Candidate_1_imm;
  wire       [3:0]    alu0Candidate_1_uop_aluOp;
  wire       [1:0]    alu0Candidate_1_uop_bruOp;
  wire       [1:0]    alu0Candidate_1_uop_cruOp;
  wire       [2:0]    alu0Candidate_1_roop_aluROOp;
  wire                alu0Candidate_1_srcReady_0;
  wire                alu0Candidate_1_srcReady_1;
  wire       [4:0]    alu1Candidate_0_robIdx;
  wire       [31:0]   alu1Candidate_0_branchInfo_predictPC;
  wire                alu1Candidate_0_branchInfo_predictResult;
  wire                alu1Candidate_0_exceptionInfo_exception;
  wire       [5:0]    alu1Candidate_0_exceptionInfo_eCode;
  wire       [0:0]    alu1Candidate_0_exceptionInfo_eSubCode;
  wire       [31:0]   alu1Candidate_0_pc;
  wire       [5:0]    alu1Candidate_0_prd;
  wire       [5:0]    alu1Candidate_0_psrc_0;
  wire       [5:0]    alu1Candidate_0_psrc_1;
  wire       [31:0]   alu1Candidate_0_imm;
  wire       [3:0]    alu1Candidate_0_uop_aluOp;
  wire       [1:0]    alu1Candidate_0_uop_bruOp;
  wire       [2:0]    alu1Candidate_0_roop_aluROOp;
  wire       [1:0]    alu1Candidate_0_roop_cruROOp;
  wire                alu1Candidate_0_srcReady_0;
  wire                alu1Candidate_0_srcReady_1;
  wire       [4:0]    alu1Candidate_1_robIdx;
  wire       [31:0]   alu1Candidate_1_branchInfo_predictPC;
  wire                alu1Candidate_1_branchInfo_predictResult;
  wire                alu1Candidate_1_exceptionInfo_exception;
  wire       [5:0]    alu1Candidate_1_exceptionInfo_eCode;
  wire       [0:0]    alu1Candidate_1_exceptionInfo_eSubCode;
  wire       [31:0]   alu1Candidate_1_pc;
  wire       [5:0]    alu1Candidate_1_prd;
  wire       [5:0]    alu1Candidate_1_psrc_0;
  wire       [5:0]    alu1Candidate_1_psrc_1;
  wire       [31:0]   alu1Candidate_1_imm;
  wire       [3:0]    alu1Candidate_1_uop_aluOp;
  wire       [1:0]    alu1Candidate_1_uop_bruOp;
  wire       [2:0]    alu1Candidate_1_roop_aluROOp;
  wire       [1:0]    alu1Candidate_1_roop_cruROOp;
  wire                alu1Candidate_1_srcReady_0;
  wire                alu1Candidate_1_srcReady_1;
  wire       [4:0]    muluCandidate_0_robIdx;
  wire       [31:0]   muluCandidate_0_branchResult_targetPC;
  wire                muluCandidate_0_branchResult_branchResult;
  wire                muluCandidate_0_branchResult_predictFail;
  wire                muluCandidate_0_exceptionInfo_exception;
  wire       [5:0]    muluCandidate_0_exceptionInfo_eCode;
  wire       [0:0]    muluCandidate_0_exceptionInfo_eSubCode;
  wire       [31:0]   muluCandidate_0_pc;
  wire       [5:0]    muluCandidate_0_prd;
  wire       [5:0]    muluCandidate_0_psrc_0;
  wire       [5:0]    muluCandidate_0_psrc_1;
  wire       [31:0]   muluCandidate_0_imm;
  wire       [1:0]    muluCandidate_0_uop_muluOp;
  wire                muluCandidate_0_srcReady_0;
  wire                muluCandidate_0_srcReady_1;
  wire       [4:0]    muluCandidate_1_robIdx;
  wire       [31:0]   muluCandidate_1_branchResult_targetPC;
  wire                muluCandidate_1_branchResult_branchResult;
  wire                muluCandidate_1_branchResult_predictFail;
  wire                muluCandidate_1_exceptionInfo_exception;
  wire       [5:0]    muluCandidate_1_exceptionInfo_eCode;
  wire       [0:0]    muluCandidate_1_exceptionInfo_eSubCode;
  wire       [31:0]   muluCandidate_1_pc;
  wire       [5:0]    muluCandidate_1_prd;
  wire       [5:0]    muluCandidate_1_psrc_0;
  wire       [5:0]    muluCandidate_1_psrc_1;
  wire       [31:0]   muluCandidate_1_imm;
  wire       [1:0]    muluCandidate_1_uop_muluOp;
  wire                muluCandidate_1_srcReady_0;
  wire                muluCandidate_1_srcReady_1;
  wire       [4:0]    divuCandidate_0_robIdx;
  wire       [31:0]   divuCandidate_0_branchResult_targetPC;
  wire                divuCandidate_0_branchResult_branchResult;
  wire                divuCandidate_0_branchResult_predictFail;
  wire                divuCandidate_0_exceptionInfo_exception;
  wire       [5:0]    divuCandidate_0_exceptionInfo_eCode;
  wire       [0:0]    divuCandidate_0_exceptionInfo_eSubCode;
  wire       [31:0]   divuCandidate_0_pc;
  wire       [5:0]    divuCandidate_0_prd;
  wire       [5:0]    divuCandidate_0_psrc_0;
  wire       [5:0]    divuCandidate_0_psrc_1;
  wire       [31:0]   divuCandidate_0_imm;
  wire       [1:0]    divuCandidate_0_uop_divuOp;
  wire                divuCandidate_0_srcReady_0;
  wire                divuCandidate_0_srcReady_1;
  wire       [4:0]    divuCandidate_1_robIdx;
  wire       [31:0]   divuCandidate_1_branchResult_targetPC;
  wire                divuCandidate_1_branchResult_branchResult;
  wire                divuCandidate_1_branchResult_predictFail;
  wire                divuCandidate_1_exceptionInfo_exception;
  wire       [5:0]    divuCandidate_1_exceptionInfo_eCode;
  wire       [0:0]    divuCandidate_1_exceptionInfo_eSubCode;
  wire       [31:0]   divuCandidate_1_pc;
  wire       [5:0]    divuCandidate_1_prd;
  wire       [5:0]    divuCandidate_1_psrc_0;
  wire       [5:0]    divuCandidate_1_psrc_1;
  wire       [31:0]   divuCandidate_1_imm;
  wire       [1:0]    divuCandidate_1_uop_divuOp;
  wire                divuCandidate_1_srcReady_0;
  wire                divuCandidate_1_srcReady_1;
  wire       [4:0]    lsuCandidate_0_robIdx;
  wire       [31:0]   lsuCandidate_0_branchResult_targetPC;
  wire                lsuCandidate_0_branchResult_branchResult;
  wire                lsuCandidate_0_branchResult_predictFail;
  wire                lsuCandidate_0_exceptionInfo_exception;
  wire       [5:0]    lsuCandidate_0_exceptionInfo_eCode;
  wire       [0:0]    lsuCandidate_0_exceptionInfo_eSubCode;
  wire       [31:0]   lsuCandidate_0_pc;
  wire       [5:0]    lsuCandidate_0_prd;
  wire       [5:0]    lsuCandidate_0_psrc_0;
  wire       [5:0]    lsuCandidate_0_psrc_1;
  wire       [31:0]   lsuCandidate_0_imm;
  wire       [3:0]    lsuCandidate_0_uop_lsuOp;
  wire       [4:0]    lsuCandidate_0_uop_lsuCoOp;
  wire       [0:0]    lsuCandidate_0_roop_lsuROOp;
  wire                lsuCandidate_0_srcReady_0;
  wire                lsuCandidate_0_srcReady_1;
  wire       [4:0]    lsuCandidate_1_robIdx;
  wire       [31:0]   lsuCandidate_1_branchResult_targetPC;
  wire                lsuCandidate_1_branchResult_branchResult;
  wire                lsuCandidate_1_branchResult_predictFail;
  wire                lsuCandidate_1_exceptionInfo_exception;
  wire       [5:0]    lsuCandidate_1_exceptionInfo_eCode;
  wire       [0:0]    lsuCandidate_1_exceptionInfo_eSubCode;
  wire       [31:0]   lsuCandidate_1_pc;
  wire       [5:0]    lsuCandidate_1_prd;
  wire       [5:0]    lsuCandidate_1_psrc_0;
  wire       [5:0]    lsuCandidate_1_psrc_1;
  wire       [31:0]   lsuCandidate_1_imm;
  wire       [3:0]    lsuCandidate_1_uop_lsuOp;
  wire       [4:0]    lsuCandidate_1_uop_lsuCoOp;
  wire       [0:0]    lsuCandidate_1_roop_lsuROOp;
  wire                lsuCandidate_1_srcReady_0;
  wire                lsuCandidate_1_srcReady_1;
  wire       [5:0]    actualSrc_0_0;
  wire       [5:0]    actualSrc_0_1;
  wire       [5:0]    actualSrc_1_0;
  wire       [5:0]    actualSrc_1_1;
  wire       [5:0]    actualRd_0;
  wire       [5:0]    actualRd_1;
  wire       [5:0]    actualpRd_0;
  wire       [5:0]    actualpRd_1;
  wire                actualSrcReady_0_0;
  wire                actualSrcReady_0_1;
  wire                actualSrcReady_1_0;
  wire                actualSrcReady_1_1;
  reg        [1:0]    _zz_actualSrcReady_1_0;
  wire       [1:0]    _zz_actualSrc_1_0;
  reg        [1:0]    _zz_actualSrc_1_0_1;
  wire       [1:0]    _zz_actualSrc_1_0_2;
  reg        [1:0]    _zz_actualSrc_1_0_3;
  reg        [1:0]    _zz_actualSrcReady_1_1;
  wire       [1:0]    _zz_actualSrc_1_1;
  reg        [1:0]    _zz_actualSrc_1_1_1;
  wire       [1:0]    _zz_actualSrc_1_1_2;
  reg        [1:0]    _zz_actualSrc_1_1_3;
  reg        [1:0]    _zz_actualpRd_1;
  wire       [1:0]    _zz_actualpRd_1_1;
  reg        [1:0]    _zz_actualpRd_1_2;
  wire       [1:0]    _zz_actualpRd_1_3;
  reg        [1:0]    _zz_actualpRd_1_4;
  wire                _zz_io_alu0IQ_payload_robIdx;
  wire       [3:0]    _zz_io_alu0IQ_payload_uop_aluOp;
  wire       [1:0]    _zz_io_alu0IQ_payload_uop_bruOp;
  wire       [1:0]    _zz_io_alu0IQ_payload_uop_cruOp;
  wire       [2:0]    _zz_io_alu0IQ_payload_roop_aluROOp;
  wire                _zz_io_alu1IQ_payload_robIdx;
  wire       [3:0]    _zz_io_alu1IQ_payload_uop_aluOp;
  wire       [1:0]    _zz_io_alu1IQ_payload_uop_bruOp;
  wire       [2:0]    _zz_io_alu1IQ_payload_roop_aluROOp;
  wire       [1:0]    _zz_io_alu1IQ_payload_roop_cruROOp;
  wire                _zz_io_muluIQ_payload_robIdx;
  wire       [1:0]    _zz_io_muluIQ_payload_uop_muluOp;
  wire                _zz_io_divuIQ_payload_robIdx;
  wire       [1:0]    _zz_io_divuIQ_payload_uop_divuOp;
  wire                _zz_io_lsuIQ_payload_robIdx;
  wire       [3:0]    _zz_io_lsuIQ_payload_uop_lsuOp;
  wire       [0:0]    _zz_io_lsuIQ_payload_roop_lsuROOp;
  `ifndef SYNTHESIS
  reg [55:0] io_input_dispatchInfo_0_fuType_string;
  reg [55:0] io_input_dispatchInfo_1_fuType_string;
  reg [71:0] io_rob_specialOp_0_string;
  reg [71:0] io_rob_specialOp_1_string;
  reg [39:0] io_alu0IQ_payload_uop_aluOp_string;
  reg [39:0] io_alu0IQ_payload_uop_bruOp_string;
  reg [31:0] io_alu0IQ_payload_uop_cruOp_string;
  reg [55:0] io_alu0IQ_payload_roop_aluROOp_string;
  reg [39:0] io_alu1IQ_payload_uop_aluOp_string;
  reg [39:0] io_alu1IQ_payload_uop_bruOp_string;
  reg [55:0] io_alu1IQ_payload_roop_aluROOp_string;
  reg [15:0] io_alu1IQ_payload_roop_cruROOp_string;
  reg [47:0] io_muluIQ_payload_uop_muluOp_string;
  reg [39:0] io_divuIQ_payload_uop_divuOp_string;
  reg [55:0] io_lsuIQ_payload_uop_lsuOp_string;
  reg [47:0] io_lsuIQ_payload_roop_lsuROOp_string;
  reg [39:0] alu0Candidate_0_uop_aluOp_string;
  reg [39:0] alu0Candidate_0_uop_bruOp_string;
  reg [31:0] alu0Candidate_0_uop_cruOp_string;
  reg [55:0] alu0Candidate_0_roop_aluROOp_string;
  reg [39:0] alu0Candidate_1_uop_aluOp_string;
  reg [39:0] alu0Candidate_1_uop_bruOp_string;
  reg [31:0] alu0Candidate_1_uop_cruOp_string;
  reg [55:0] alu0Candidate_1_roop_aluROOp_string;
  reg [39:0] alu1Candidate_0_uop_aluOp_string;
  reg [39:0] alu1Candidate_0_uop_bruOp_string;
  reg [55:0] alu1Candidate_0_roop_aluROOp_string;
  reg [15:0] alu1Candidate_0_roop_cruROOp_string;
  reg [39:0] alu1Candidate_1_uop_aluOp_string;
  reg [39:0] alu1Candidate_1_uop_bruOp_string;
  reg [55:0] alu1Candidate_1_roop_aluROOp_string;
  reg [15:0] alu1Candidate_1_roop_cruROOp_string;
  reg [47:0] muluCandidate_0_uop_muluOp_string;
  reg [47:0] muluCandidate_1_uop_muluOp_string;
  reg [39:0] divuCandidate_0_uop_divuOp_string;
  reg [39:0] divuCandidate_1_uop_divuOp_string;
  reg [55:0] lsuCandidate_0_uop_lsuOp_string;
  reg [47:0] lsuCandidate_0_roop_lsuROOp_string;
  reg [55:0] lsuCandidate_1_uop_lsuOp_string;
  reg [47:0] lsuCandidate_1_roop_lsuROOp_string;
  reg [39:0] _zz_io_alu0IQ_payload_uop_aluOp_string;
  reg [39:0] _zz_io_alu0IQ_payload_uop_bruOp_string;
  reg [31:0] _zz_io_alu0IQ_payload_uop_cruOp_string;
  reg [55:0] _zz_io_alu0IQ_payload_roop_aluROOp_string;
  reg [39:0] _zz_io_alu1IQ_payload_uop_aluOp_string;
  reg [39:0] _zz_io_alu1IQ_payload_uop_bruOp_string;
  reg [55:0] _zz_io_alu1IQ_payload_roop_aluROOp_string;
  reg [15:0] _zz_io_alu1IQ_payload_roop_cruROOp_string;
  reg [47:0] _zz_io_muluIQ_payload_uop_muluOp_string;
  reg [39:0] _zz_io_divuIQ_payload_uop_divuOp_string;
  reg [55:0] _zz_io_lsuIQ_payload_uop_lsuOp_string;
  reg [47:0] _zz_io_lsuIQ_payload_roop_lsuROOp_string;
  `endif


  assign _zz_alu0Sel_1 = (_zz_alu0Sel - 2'b01);
  assign _zz_alu1Sel_1 = (_zz_alu1Sel - 2'b01);
  assign _zz_muluReq_ohFirst_masked = (muluReq_ohFirst_input - 2'b01);
  assign _zz_divuReq_ohFirst_masked = (divuReq_ohFirst_input - 2'b01);
  assign _zz_lsuReq_ohFirst_masked = (lsuReq_ohFirst_input - 2'b01);
  assign _zz__zz_actualSrc_1_0_2 = (_zz_actualSrc_1_0_1 - 2'b01);
  assign _zz__zz_actualSrc_1_1_2 = (_zz_actualSrc_1_1_1 - 2'b01);
  assign _zz__zz_actualpRd_1_3 = (_zz_actualpRd_1_2 - 2'b01);
  assign _zz_freelistRdShuffle_1_2 = needRd[0];
  assign _zz_freelistAvail_1 = needRd[0];
  assign _zz_io_freelist_disPatchNum_1 = {dispatchMask[1],dispatchMask[0]};
  Decoder decoder_0 (
    .io_info_inst                     (io_input_info_0_inst[31:0]                ), //i
    .io_info_branchInfo_predictPC     (io_input_info_0_branchInfo_predictPC[31:0]), //i
    .io_info_branchInfo_predictResult (io_input_info_0_branchInfo_predictResult  ), //i
    .io_info_exceptionInfo_exception  (io_input_info_0_exceptionInfo_exception   ), //i
    .io_info_exceptionInfo_eCode      (io_input_info_0_exceptionInfo_eCode[5:0]  ), //i
    .io_info_exceptionInfo_eSubCode   (io_input_info_0_exceptionInfo_eSubCode    ), //i
    .io_info_pc                       (io_input_info_0_pc[31:0]                  ), //i
    ._zz_when_Decoder_l40             (_zz_when_Decoder_l40[1:0]                 ), //i
    .io_branchInfo_predictPC          (decoder_0_io_branchInfo_predictPC[31:0]   ), //o
    .io_branchInfo_predictResult      (decoder_0_io_branchInfo_predictResult     ), //o
    .io_branchResult_targetPC         (decoder_0_io_branchResult_targetPC[31:0]  ), //o
    .io_branchResult_branchResult     (decoder_0_io_branchResult_branchResult    ), //o
    .io_branchResult_predictFail      (decoder_0_io_branchResult_predictFail     ), //o
    .io_exceptionInfo_exception       (decoder_0_io_exceptionInfo_exception      ), //o
    .io_exceptionInfo_eCode           (decoder_0_io_exceptionInfo_eCode[5:0]     ), //o
    .io_exceptionInfo_eSubCode        (decoder_0_io_exceptionInfo_eSubCode       ), //o
    .io_pc                            (decoder_0_io_pc[31:0]                     ), //o
    .io_specialOp                     (decoder_0_io_specialOp[3:0]               ), //o
    .io_imm                           (decoder_0_io_imm[31:0]                    ), //o
    .io_uopALU0_aluOp                 (decoder_0_io_uopALU0_aluOp[3:0]           ), //o
    .io_uopALU0_bruOp                 (decoder_0_io_uopALU0_bruOp[1:0]           ), //o
    .io_uopALU0_cruOp                 (decoder_0_io_uopALU0_cruOp[1:0]           ), //o
    .io_uopALU1_aluOp                 (decoder_0_io_uopALU1_aluOp[3:0]           ), //o
    .io_uopALU1_bruOp                 (decoder_0_io_uopALU1_bruOp[1:0]           ), //o
    .io_uopMULU_muluOp                (decoder_0_io_uopMULU_muluOp[1:0]          ), //o
    .io_uopDIVU_divuOp                (decoder_0_io_uopDIVU_divuOp[1:0]          ), //o
    .io_uopLSU_lsuOp                  (decoder_0_io_uopLSU_lsuOp[3:0]            ), //o
    .io_uopLSU_lsuCoOp                (decoder_0_io_uopLSU_lsuCoOp[4:0]          ), //o
    .io_roopALU0_aluROOp              (decoder_0_io_roopALU0_aluROOp[2:0]        ), //o
    .io_roopALU1_aluROOp              (decoder_0_io_roopALU1_aluROOp[2:0]        ), //o
    .io_roopALU1_cruROOp              (decoder_0_io_roopALU1_cruROOp[1:0]        ), //o
    .io_roopLSU_lsuROOp               (decoder_0_io_roopLSU_lsuROOp              )  //o
  );
  Decoder decoder_1_1 (
    .io_info_inst                     (io_input_info_1_inst[31:0]                ), //i
    .io_info_branchInfo_predictPC     (io_input_info_1_branchInfo_predictPC[31:0]), //i
    .io_info_branchInfo_predictResult (io_input_info_1_branchInfo_predictResult  ), //i
    .io_info_exceptionInfo_exception  (io_input_info_1_exceptionInfo_exception   ), //i
    .io_info_exceptionInfo_eCode      (io_input_info_1_exceptionInfo_eCode[5:0]  ), //i
    .io_info_exceptionInfo_eSubCode   (io_input_info_1_exceptionInfo_eSubCode    ), //i
    .io_info_pc                       (io_input_info_1_pc[31:0]                  ), //i
    ._zz_when_Decoder_l40             (_zz_when_Decoder_l40[1:0]                 ), //i
    .io_branchInfo_predictPC          (decoder_1_1_io_branchInfo_predictPC[31:0] ), //o
    .io_branchInfo_predictResult      (decoder_1_1_io_branchInfo_predictResult   ), //o
    .io_branchResult_targetPC         (decoder_1_1_io_branchResult_targetPC[31:0]), //o
    .io_branchResult_branchResult     (decoder_1_1_io_branchResult_branchResult  ), //o
    .io_branchResult_predictFail      (decoder_1_1_io_branchResult_predictFail   ), //o
    .io_exceptionInfo_exception       (decoder_1_1_io_exceptionInfo_exception    ), //o
    .io_exceptionInfo_eCode           (decoder_1_1_io_exceptionInfo_eCode[5:0]   ), //o
    .io_exceptionInfo_eSubCode        (decoder_1_1_io_exceptionInfo_eSubCode     ), //o
    .io_pc                            (decoder_1_1_io_pc[31:0]                   ), //o
    .io_specialOp                     (decoder_1_1_io_specialOp[3:0]             ), //o
    .io_imm                           (decoder_1_1_io_imm[31:0]                  ), //o
    .io_uopALU0_aluOp                 (decoder_1_1_io_uopALU0_aluOp[3:0]         ), //o
    .io_uopALU0_bruOp                 (decoder_1_1_io_uopALU0_bruOp[1:0]         ), //o
    .io_uopALU0_cruOp                 (decoder_1_1_io_uopALU0_cruOp[1:0]         ), //o
    .io_uopALU1_aluOp                 (decoder_1_1_io_uopALU1_aluOp[3:0]         ), //o
    .io_uopALU1_bruOp                 (decoder_1_1_io_uopALU1_bruOp[1:0]         ), //o
    .io_uopMULU_muluOp                (decoder_1_1_io_uopMULU_muluOp[1:0]        ), //o
    .io_uopDIVU_divuOp                (decoder_1_1_io_uopDIVU_divuOp[1:0]        ), //o
    .io_uopLSU_lsuOp                  (decoder_1_1_io_uopLSU_lsuOp[3:0]          ), //o
    .io_uopLSU_lsuCoOp                (decoder_1_1_io_uopLSU_lsuCoOp[4:0]        ), //o
    .io_roopALU0_aluROOp              (decoder_1_1_io_roopALU0_aluROOp[2:0]      ), //o
    .io_roopALU1_aluROOp              (decoder_1_1_io_roopALU1_aluROOp[2:0]      ), //o
    .io_roopALU1_cruROOp              (decoder_1_1_io_roopALU1_cruROOp[1:0]      ), //o
    .io_roopLSU_lsuROOp               (decoder_1_1_io_roopLSU_lsuROOp            )  //o
  );
  always @(*) begin
    case(_zz_freelistRdShuffle_1_1)
      1'b0 : _zz_freelistRdShuffle_1 = io_freelist_prfIdx_0;
      default : _zz_freelistRdShuffle_1 = io_freelist_prfIdx_1;
    endcase
  end

  always @(*) begin
    case(_zz_freelistRdShuffle_1_2)
      1'b0 : _zz_freelistRdShuffle_1_1 = 1'b0;
      default : _zz_freelistRdShuffle_1_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_freelistAvail_1)
      1'b0 : _zz_freelistAvail = 1'b0;
      default : _zz_freelistAvail = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_io_freelist_disPatchNum_1)
      2'b00 : _zz_io_freelist_disPatchNum = 2'b00;
      2'b01 : _zz_io_freelist_disPatchNum = 2'b01;
      2'b10 : _zz_io_freelist_disPatchNum = 2'b01;
      default : _zz_io_freelist_disPatchNum = 2'b10;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_dispatchInfo_0_fuType)
      FUType_alu : io_input_dispatchInfo_0_fuType_string = "alu    ";
      FUType_csr : io_input_dispatchInfo_0_fuType_string = "csr    ";
      FUType_counter : io_input_dispatchInfo_0_fuType_string = "counter";
      FUType_lsu : io_input_dispatchInfo_0_fuType_string = "lsu    ";
      FUType_mulu : io_input_dispatchInfo_0_fuType_string = "mulu   ";
      FUType_divu : io_input_dispatchInfo_0_fuType_string = "divu   ";
      default : io_input_dispatchInfo_0_fuType_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_input_dispatchInfo_1_fuType)
      FUType_alu : io_input_dispatchInfo_1_fuType_string = "alu    ";
      FUType_csr : io_input_dispatchInfo_1_fuType_string = "csr    ";
      FUType_counter : io_input_dispatchInfo_1_fuType_string = "counter";
      FUType_lsu : io_input_dispatchInfo_1_fuType_string = "lsu    ";
      FUType_mulu : io_input_dispatchInfo_1_fuType_string = "mulu   ";
      FUType_divu : io_input_dispatchInfo_1_fuType_string = "divu   ";
      default : io_input_dispatchInfo_1_fuType_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_rob_specialOp_0)
      ROBSpecialOp_nop : io_rob_specialOp_0_string = "nop      ";
      ROBSpecialOp_bpuUpdate : io_rob_specialOp_0_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : io_rob_specialOp_0_string = "lsuAction";
      ROBSpecialOp_ll : io_rob_specialOp_0_string = "ll       ";
      ROBSpecialOp_writeCSR : io_rob_specialOp_0_string = "writeCSR ";
      ROBSpecialOp_ertn : io_rob_specialOp_0_string = "ertn     ";
      ROBSpecialOp_idle : io_rob_specialOp_0_string = "idle     ";
      ROBSpecialOp_readCSR : io_rob_specialOp_0_string = "readCSR  ";
      ROBSpecialOp_readCNT : io_rob_specialOp_0_string = "readCNT  ";
      default : io_rob_specialOp_0_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_rob_specialOp_1)
      ROBSpecialOp_nop : io_rob_specialOp_1_string = "nop      ";
      ROBSpecialOp_bpuUpdate : io_rob_specialOp_1_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : io_rob_specialOp_1_string = "lsuAction";
      ROBSpecialOp_ll : io_rob_specialOp_1_string = "ll       ";
      ROBSpecialOp_writeCSR : io_rob_specialOp_1_string = "writeCSR ";
      ROBSpecialOp_ertn : io_rob_specialOp_1_string = "ertn     ";
      ROBSpecialOp_idle : io_rob_specialOp_1_string = "idle     ";
      ROBSpecialOp_readCSR : io_rob_specialOp_1_string = "readCSR  ";
      ROBSpecialOp_readCNT : io_rob_specialOp_1_string = "readCNT  ";
      default : io_rob_specialOp_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_alu0IQ_payload_uop_aluOp)
      ALUOp_add : io_alu0IQ_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_alu0IQ_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_alu0IQ_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_alu0IQ_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_alu0IQ_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_alu0IQ_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_alu0IQ_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_alu0IQ_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_alu0IQ_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_alu0IQ_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_alu0IQ_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_alu0IQ_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_alu0IQ_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_alu0IQ_payload_uop_aluOp_string = "passb";
      default : io_alu0IQ_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_alu0IQ_payload_uop_bruOp)
      BRUOp_nop : io_alu0IQ_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_alu0IQ_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_alu0IQ_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_alu0IQ_payload_uop_bruOp_string = "ncadd";
      default : io_alu0IQ_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_alu0IQ_payload_uop_cruOp)
      CRUOp_nop : io_alu0IQ_payload_uop_cruOp_string = "nop ";
      CRUOp_pass : io_alu0IQ_payload_uop_cruOp_string = "pass";
      CRUOp_mask : io_alu0IQ_payload_uop_cruOp_string = "mask";
      default : io_alu0IQ_payload_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(io_alu0IQ_payload_roop_aluROOp)
      ALUROOp_reg_1 : io_alu0IQ_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : io_alu0IQ_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : io_alu0IQ_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : io_alu0IQ_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : io_alu0IQ_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : io_alu0IQ_payload_roop_aluROOp_string = "linkreg";
      default : io_alu0IQ_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_alu1IQ_payload_uop_aluOp)
      ALUOp_add : io_alu1IQ_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : io_alu1IQ_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : io_alu1IQ_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : io_alu1IQ_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : io_alu1IQ_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_alu1IQ_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : io_alu1IQ_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : io_alu1IQ_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_alu1IQ_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_alu1IQ_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_alu1IQ_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_alu1IQ_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : io_alu1IQ_payload_uop_aluOp_string = "passa";
      ALUOp_passb : io_alu1IQ_payload_uop_aluOp_string = "passb";
      default : io_alu1IQ_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_alu1IQ_payload_uop_bruOp)
      BRUOp_nop : io_alu1IQ_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : io_alu1IQ_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : io_alu1IQ_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : io_alu1IQ_payload_uop_bruOp_string = "ncadd";
      default : io_alu1IQ_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_alu1IQ_payload_roop_aluROOp)
      ALUROOp_reg_1 : io_alu1IQ_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : io_alu1IQ_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : io_alu1IQ_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : io_alu1IQ_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : io_alu1IQ_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : io_alu1IQ_payload_roop_aluROOp_string = "linkreg";
      default : io_alu1IQ_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_alu1IQ_payload_roop_cruROOp)
      CRUROOp_id : io_alu1IQ_payload_roop_cruROOp_string = "id";
      CRUROOp_lo : io_alu1IQ_payload_roop_cruROOp_string = "lo";
      CRUROOp_hi : io_alu1IQ_payload_roop_cruROOp_string = "hi";
      default : io_alu1IQ_payload_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(io_muluIQ_payload_uop_muluOp)
      MULUOp_mullo : io_muluIQ_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : io_muluIQ_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : io_muluIQ_payload_uop_muluOp_string = "mulhiu";
      default : io_muluIQ_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_divuIQ_payload_uop_divuOp)
      DIVUOp_div : io_divuIQ_payload_uop_divuOp_string = "div  ";
      DIVUOp_divu : io_divuIQ_payload_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : io_divuIQ_payload_uop_divuOp_string = "mod_1";
      DIVUOp_modu : io_divuIQ_payload_uop_divuOp_string = "modu ";
      default : io_divuIQ_payload_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_lsuIQ_payload_uop_lsuOp)
      LSUOp_cacop : io_lsuIQ_payload_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : io_lsuIQ_payload_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : io_lsuIQ_payload_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : io_lsuIQ_payload_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : io_lsuIQ_payload_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : io_lsuIQ_payload_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : io_lsuIQ_payload_uop_lsuOp_string = "ll     ";
      LSUOp_sc : io_lsuIQ_payload_uop_lsuOp_string = "sc     ";
      LSUOp_ld : io_lsuIQ_payload_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : io_lsuIQ_payload_uop_lsuOp_string = "ldu    ";
      LSUOp_st : io_lsuIQ_payload_uop_lsuOp_string = "st     ";
      LSUOp_preld : io_lsuIQ_payload_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : io_lsuIQ_payload_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : io_lsuIQ_payload_uop_lsuOp_string = "ibar   ";
      default : io_lsuIQ_payload_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_lsuIQ_payload_roop_lsuROOp)
      LSUROOp_reg_1 : io_lsuIQ_payload_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : io_lsuIQ_payload_roop_lsuROOp_string = "regimm";
      default : io_lsuIQ_payload_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(alu0Candidate_0_uop_aluOp)
      ALUOp_add : alu0Candidate_0_uop_aluOp_string = "add  ";
      ALUOp_sub : alu0Candidate_0_uop_aluOp_string = "sub  ";
      ALUOp_slt : alu0Candidate_0_uop_aluOp_string = "slt  ";
      ALUOp_sltu : alu0Candidate_0_uop_aluOp_string = "sltu ";
      ALUOp_eq : alu0Candidate_0_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : alu0Candidate_0_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : alu0Candidate_0_uop_aluOp_string = "and_1";
      ALUOp_or_1 : alu0Candidate_0_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : alu0Candidate_0_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : alu0Candidate_0_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : alu0Candidate_0_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : alu0Candidate_0_uop_aluOp_string = "sra_1";
      ALUOp_passa : alu0Candidate_0_uop_aluOp_string = "passa";
      ALUOp_passb : alu0Candidate_0_uop_aluOp_string = "passb";
      default : alu0Candidate_0_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(alu0Candidate_0_uop_bruOp)
      BRUOp_nop : alu0Candidate_0_uop_bruOp_string = "nop  ";
      BRUOp_add : alu0Candidate_0_uop_bruOp_string = "add  ";
      BRUOp_cadd : alu0Candidate_0_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : alu0Candidate_0_uop_bruOp_string = "ncadd";
      default : alu0Candidate_0_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(alu0Candidate_0_uop_cruOp)
      CRUOp_nop : alu0Candidate_0_uop_cruOp_string = "nop ";
      CRUOp_pass : alu0Candidate_0_uop_cruOp_string = "pass";
      CRUOp_mask : alu0Candidate_0_uop_cruOp_string = "mask";
      default : alu0Candidate_0_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(alu0Candidate_0_roop_aluROOp)
      ALUROOp_reg_1 : alu0Candidate_0_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : alu0Candidate_0_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : alu0Candidate_0_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : alu0Candidate_0_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : alu0Candidate_0_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : alu0Candidate_0_roop_aluROOp_string = "linkreg";
      default : alu0Candidate_0_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(alu0Candidate_1_uop_aluOp)
      ALUOp_add : alu0Candidate_1_uop_aluOp_string = "add  ";
      ALUOp_sub : alu0Candidate_1_uop_aluOp_string = "sub  ";
      ALUOp_slt : alu0Candidate_1_uop_aluOp_string = "slt  ";
      ALUOp_sltu : alu0Candidate_1_uop_aluOp_string = "sltu ";
      ALUOp_eq : alu0Candidate_1_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : alu0Candidate_1_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : alu0Candidate_1_uop_aluOp_string = "and_1";
      ALUOp_or_1 : alu0Candidate_1_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : alu0Candidate_1_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : alu0Candidate_1_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : alu0Candidate_1_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : alu0Candidate_1_uop_aluOp_string = "sra_1";
      ALUOp_passa : alu0Candidate_1_uop_aluOp_string = "passa";
      ALUOp_passb : alu0Candidate_1_uop_aluOp_string = "passb";
      default : alu0Candidate_1_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(alu0Candidate_1_uop_bruOp)
      BRUOp_nop : alu0Candidate_1_uop_bruOp_string = "nop  ";
      BRUOp_add : alu0Candidate_1_uop_bruOp_string = "add  ";
      BRUOp_cadd : alu0Candidate_1_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : alu0Candidate_1_uop_bruOp_string = "ncadd";
      default : alu0Candidate_1_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(alu0Candidate_1_uop_cruOp)
      CRUOp_nop : alu0Candidate_1_uop_cruOp_string = "nop ";
      CRUOp_pass : alu0Candidate_1_uop_cruOp_string = "pass";
      CRUOp_mask : alu0Candidate_1_uop_cruOp_string = "mask";
      default : alu0Candidate_1_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(alu0Candidate_1_roop_aluROOp)
      ALUROOp_reg_1 : alu0Candidate_1_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : alu0Candidate_1_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : alu0Candidate_1_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : alu0Candidate_1_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : alu0Candidate_1_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : alu0Candidate_1_roop_aluROOp_string = "linkreg";
      default : alu0Candidate_1_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(alu1Candidate_0_uop_aluOp)
      ALUOp_add : alu1Candidate_0_uop_aluOp_string = "add  ";
      ALUOp_sub : alu1Candidate_0_uop_aluOp_string = "sub  ";
      ALUOp_slt : alu1Candidate_0_uop_aluOp_string = "slt  ";
      ALUOp_sltu : alu1Candidate_0_uop_aluOp_string = "sltu ";
      ALUOp_eq : alu1Candidate_0_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : alu1Candidate_0_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : alu1Candidate_0_uop_aluOp_string = "and_1";
      ALUOp_or_1 : alu1Candidate_0_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : alu1Candidate_0_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : alu1Candidate_0_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : alu1Candidate_0_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : alu1Candidate_0_uop_aluOp_string = "sra_1";
      ALUOp_passa : alu1Candidate_0_uop_aluOp_string = "passa";
      ALUOp_passb : alu1Candidate_0_uop_aluOp_string = "passb";
      default : alu1Candidate_0_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(alu1Candidate_0_uop_bruOp)
      BRUOp_nop : alu1Candidate_0_uop_bruOp_string = "nop  ";
      BRUOp_add : alu1Candidate_0_uop_bruOp_string = "add  ";
      BRUOp_cadd : alu1Candidate_0_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : alu1Candidate_0_uop_bruOp_string = "ncadd";
      default : alu1Candidate_0_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(alu1Candidate_0_roop_aluROOp)
      ALUROOp_reg_1 : alu1Candidate_0_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : alu1Candidate_0_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : alu1Candidate_0_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : alu1Candidate_0_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : alu1Candidate_0_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : alu1Candidate_0_roop_aluROOp_string = "linkreg";
      default : alu1Candidate_0_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(alu1Candidate_0_roop_cruROOp)
      CRUROOp_id : alu1Candidate_0_roop_cruROOp_string = "id";
      CRUROOp_lo : alu1Candidate_0_roop_cruROOp_string = "lo";
      CRUROOp_hi : alu1Candidate_0_roop_cruROOp_string = "hi";
      default : alu1Candidate_0_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(alu1Candidate_1_uop_aluOp)
      ALUOp_add : alu1Candidate_1_uop_aluOp_string = "add  ";
      ALUOp_sub : alu1Candidate_1_uop_aluOp_string = "sub  ";
      ALUOp_slt : alu1Candidate_1_uop_aluOp_string = "slt  ";
      ALUOp_sltu : alu1Candidate_1_uop_aluOp_string = "sltu ";
      ALUOp_eq : alu1Candidate_1_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : alu1Candidate_1_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : alu1Candidate_1_uop_aluOp_string = "and_1";
      ALUOp_or_1 : alu1Candidate_1_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : alu1Candidate_1_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : alu1Candidate_1_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : alu1Candidate_1_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : alu1Candidate_1_uop_aluOp_string = "sra_1";
      ALUOp_passa : alu1Candidate_1_uop_aluOp_string = "passa";
      ALUOp_passb : alu1Candidate_1_uop_aluOp_string = "passb";
      default : alu1Candidate_1_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(alu1Candidate_1_uop_bruOp)
      BRUOp_nop : alu1Candidate_1_uop_bruOp_string = "nop  ";
      BRUOp_add : alu1Candidate_1_uop_bruOp_string = "add  ";
      BRUOp_cadd : alu1Candidate_1_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : alu1Candidate_1_uop_bruOp_string = "ncadd";
      default : alu1Candidate_1_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(alu1Candidate_1_roop_aluROOp)
      ALUROOp_reg_1 : alu1Candidate_1_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : alu1Candidate_1_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : alu1Candidate_1_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : alu1Candidate_1_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : alu1Candidate_1_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : alu1Candidate_1_roop_aluROOp_string = "linkreg";
      default : alu1Candidate_1_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(alu1Candidate_1_roop_cruROOp)
      CRUROOp_id : alu1Candidate_1_roop_cruROOp_string = "id";
      CRUROOp_lo : alu1Candidate_1_roop_cruROOp_string = "lo";
      CRUROOp_hi : alu1Candidate_1_roop_cruROOp_string = "hi";
      default : alu1Candidate_1_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(muluCandidate_0_uop_muluOp)
      MULUOp_mullo : muluCandidate_0_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : muluCandidate_0_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : muluCandidate_0_uop_muluOp_string = "mulhiu";
      default : muluCandidate_0_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(muluCandidate_1_uop_muluOp)
      MULUOp_mullo : muluCandidate_1_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : muluCandidate_1_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : muluCandidate_1_uop_muluOp_string = "mulhiu";
      default : muluCandidate_1_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(divuCandidate_0_uop_divuOp)
      DIVUOp_div : divuCandidate_0_uop_divuOp_string = "div  ";
      DIVUOp_divu : divuCandidate_0_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : divuCandidate_0_uop_divuOp_string = "mod_1";
      DIVUOp_modu : divuCandidate_0_uop_divuOp_string = "modu ";
      default : divuCandidate_0_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(divuCandidate_1_uop_divuOp)
      DIVUOp_div : divuCandidate_1_uop_divuOp_string = "div  ";
      DIVUOp_divu : divuCandidate_1_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : divuCandidate_1_uop_divuOp_string = "mod_1";
      DIVUOp_modu : divuCandidate_1_uop_divuOp_string = "modu ";
      default : divuCandidate_1_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(lsuCandidate_0_uop_lsuOp)
      LSUOp_cacop : lsuCandidate_0_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : lsuCandidate_0_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : lsuCandidate_0_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : lsuCandidate_0_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : lsuCandidate_0_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : lsuCandidate_0_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : lsuCandidate_0_uop_lsuOp_string = "ll     ";
      LSUOp_sc : lsuCandidate_0_uop_lsuOp_string = "sc     ";
      LSUOp_ld : lsuCandidate_0_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : lsuCandidate_0_uop_lsuOp_string = "ldu    ";
      LSUOp_st : lsuCandidate_0_uop_lsuOp_string = "st     ";
      LSUOp_preld : lsuCandidate_0_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : lsuCandidate_0_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : lsuCandidate_0_uop_lsuOp_string = "ibar   ";
      default : lsuCandidate_0_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(lsuCandidate_0_roop_lsuROOp)
      LSUROOp_reg_1 : lsuCandidate_0_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : lsuCandidate_0_roop_lsuROOp_string = "regimm";
      default : lsuCandidate_0_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(lsuCandidate_1_uop_lsuOp)
      LSUOp_cacop : lsuCandidate_1_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : lsuCandidate_1_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : lsuCandidate_1_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : lsuCandidate_1_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : lsuCandidate_1_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : lsuCandidate_1_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : lsuCandidate_1_uop_lsuOp_string = "ll     ";
      LSUOp_sc : lsuCandidate_1_uop_lsuOp_string = "sc     ";
      LSUOp_ld : lsuCandidate_1_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : lsuCandidate_1_uop_lsuOp_string = "ldu    ";
      LSUOp_st : lsuCandidate_1_uop_lsuOp_string = "st     ";
      LSUOp_preld : lsuCandidate_1_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : lsuCandidate_1_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : lsuCandidate_1_uop_lsuOp_string = "ibar   ";
      default : lsuCandidate_1_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(lsuCandidate_1_roop_lsuROOp)
      LSUROOp_reg_1 : lsuCandidate_1_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : lsuCandidate_1_roop_lsuROOp_string = "regimm";
      default : lsuCandidate_1_roop_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_alu0IQ_payload_uop_aluOp)
      ALUOp_add : _zz_io_alu0IQ_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : _zz_io_alu0IQ_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : _zz_io_alu0IQ_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : _zz_io_alu0IQ_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : _zz_io_alu0IQ_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : _zz_io_alu0IQ_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : _zz_io_alu0IQ_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : _zz_io_alu0IQ_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : _zz_io_alu0IQ_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : _zz_io_alu0IQ_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : _zz_io_alu0IQ_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : _zz_io_alu0IQ_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : _zz_io_alu0IQ_payload_uop_aluOp_string = "passa";
      ALUOp_passb : _zz_io_alu0IQ_payload_uop_aluOp_string = "passb";
      default : _zz_io_alu0IQ_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_alu0IQ_payload_uop_bruOp)
      BRUOp_nop : _zz_io_alu0IQ_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : _zz_io_alu0IQ_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : _zz_io_alu0IQ_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : _zz_io_alu0IQ_payload_uop_bruOp_string = "ncadd";
      default : _zz_io_alu0IQ_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_alu0IQ_payload_uop_cruOp)
      CRUOp_nop : _zz_io_alu0IQ_payload_uop_cruOp_string = "nop ";
      CRUOp_pass : _zz_io_alu0IQ_payload_uop_cruOp_string = "pass";
      CRUOp_mask : _zz_io_alu0IQ_payload_uop_cruOp_string = "mask";
      default : _zz_io_alu0IQ_payload_uop_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_io_alu0IQ_payload_roop_aluROOp)
      ALUROOp_reg_1 : _zz_io_alu0IQ_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : _zz_io_alu0IQ_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : _zz_io_alu0IQ_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : _zz_io_alu0IQ_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : _zz_io_alu0IQ_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : _zz_io_alu0IQ_payload_roop_aluROOp_string = "linkreg";
      default : _zz_io_alu0IQ_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(_zz_io_alu1IQ_payload_uop_aluOp)
      ALUOp_add : _zz_io_alu1IQ_payload_uop_aluOp_string = "add  ";
      ALUOp_sub : _zz_io_alu1IQ_payload_uop_aluOp_string = "sub  ";
      ALUOp_slt : _zz_io_alu1IQ_payload_uop_aluOp_string = "slt  ";
      ALUOp_sltu : _zz_io_alu1IQ_payload_uop_aluOp_string = "sltu ";
      ALUOp_eq : _zz_io_alu1IQ_payload_uop_aluOp_string = "eq   ";
      ALUOp_nor_1 : _zz_io_alu1IQ_payload_uop_aluOp_string = "nor_1";
      ALUOp_and_1 : _zz_io_alu1IQ_payload_uop_aluOp_string = "and_1";
      ALUOp_or_1 : _zz_io_alu1IQ_payload_uop_aluOp_string = "or_1 ";
      ALUOp_xor_1 : _zz_io_alu1IQ_payload_uop_aluOp_string = "xor_1";
      ALUOp_sll_1 : _zz_io_alu1IQ_payload_uop_aluOp_string = "sll_1";
      ALUOp_srl_1 : _zz_io_alu1IQ_payload_uop_aluOp_string = "srl_1";
      ALUOp_sra_1 : _zz_io_alu1IQ_payload_uop_aluOp_string = "sra_1";
      ALUOp_passa : _zz_io_alu1IQ_payload_uop_aluOp_string = "passa";
      ALUOp_passb : _zz_io_alu1IQ_payload_uop_aluOp_string = "passb";
      default : _zz_io_alu1IQ_payload_uop_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_alu1IQ_payload_uop_bruOp)
      BRUOp_nop : _zz_io_alu1IQ_payload_uop_bruOp_string = "nop  ";
      BRUOp_add : _zz_io_alu1IQ_payload_uop_bruOp_string = "add  ";
      BRUOp_cadd : _zz_io_alu1IQ_payload_uop_bruOp_string = "cadd ";
      BRUOp_ncadd : _zz_io_alu1IQ_payload_uop_bruOp_string = "ncadd";
      default : _zz_io_alu1IQ_payload_uop_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_alu1IQ_payload_roop_aluROOp)
      ALUROOp_reg_1 : _zz_io_alu1IQ_payload_roop_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : _zz_io_alu1IQ_payload_roop_aluROOp_string = "regimm ";
      ALUROOp_pcimm : _zz_io_alu1IQ_payload_roop_aluROOp_string = "pcimm  ";
      ALUROOp_csr : _zz_io_alu1IQ_payload_roop_aluROOp_string = "csr    ";
      ALUROOp_linkpc : _zz_io_alu1IQ_payload_roop_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : _zz_io_alu1IQ_payload_roop_aluROOp_string = "linkreg";
      default : _zz_io_alu1IQ_payload_roop_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(_zz_io_alu1IQ_payload_roop_cruROOp)
      CRUROOp_id : _zz_io_alu1IQ_payload_roop_cruROOp_string = "id";
      CRUROOp_lo : _zz_io_alu1IQ_payload_roop_cruROOp_string = "lo";
      CRUROOp_hi : _zz_io_alu1IQ_payload_roop_cruROOp_string = "hi";
      default : _zz_io_alu1IQ_payload_roop_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(_zz_io_muluIQ_payload_uop_muluOp)
      MULUOp_mullo : _zz_io_muluIQ_payload_uop_muluOp_string = "mullo ";
      MULUOp_mulhi : _zz_io_muluIQ_payload_uop_muluOp_string = "mulhi ";
      MULUOp_mulhiu : _zz_io_muluIQ_payload_uop_muluOp_string = "mulhiu";
      default : _zz_io_muluIQ_payload_uop_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_divuIQ_payload_uop_divuOp)
      DIVUOp_div : _zz_io_divuIQ_payload_uop_divuOp_string = "div  ";
      DIVUOp_divu : _zz_io_divuIQ_payload_uop_divuOp_string = "divu ";
      DIVUOp_mod_1 : _zz_io_divuIQ_payload_uop_divuOp_string = "mod_1";
      DIVUOp_modu : _zz_io_divuIQ_payload_uop_divuOp_string = "modu ";
      default : _zz_io_divuIQ_payload_uop_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_io_lsuIQ_payload_uop_lsuOp)
      LSUOp_cacop : _zz_io_lsuIQ_payload_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : _zz_io_lsuIQ_payload_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : _zz_io_lsuIQ_payload_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : _zz_io_lsuIQ_payload_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : _zz_io_lsuIQ_payload_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : _zz_io_lsuIQ_payload_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : _zz_io_lsuIQ_payload_uop_lsuOp_string = "ll     ";
      LSUOp_sc : _zz_io_lsuIQ_payload_uop_lsuOp_string = "sc     ";
      LSUOp_ld : _zz_io_lsuIQ_payload_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : _zz_io_lsuIQ_payload_uop_lsuOp_string = "ldu    ";
      LSUOp_st : _zz_io_lsuIQ_payload_uop_lsuOp_string = "st     ";
      LSUOp_preld : _zz_io_lsuIQ_payload_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : _zz_io_lsuIQ_payload_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : _zz_io_lsuIQ_payload_uop_lsuOp_string = "ibar   ";
      default : _zz_io_lsuIQ_payload_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(_zz_io_lsuIQ_payload_roop_lsuROOp)
      LSUROOp_reg_1 : _zz_io_lsuIQ_payload_roop_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : _zz_io_lsuIQ_payload_roop_lsuROOp_string = "regimm";
      default : _zz_io_lsuIQ_payload_roop_lsuROOp_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    needRd[0] = (io_input_dispatchInfo_0_ard != 5'h00);
    needRd[1] = (io_input_dispatchInfo_1_ard != 5'h00);
  end

  assign when_Dispatcher_l34 = needRd[0];
  always @(*) begin
    if(when_Dispatcher_l34) begin
      freelistRdShuffle_0 = io_freelist_prfIdx_0;
    end else begin
      freelistRdShuffle_0 = 6'h00;
    end
  end

  always @(*) begin
    if(when_Dispatcher_l34) begin
      freelistAvail[0] = io_freelist_availMask[0];
    end else begin
      freelistAvail[0] = 1'b1;
    end
    if(when_Dispatcher_l42) begin
      freelistAvail[1] = io_freelist_availMask[_zz_freelistAvail];
    end else begin
      freelistAvail[1] = 1'b1;
    end
  end

  assign when_Dispatcher_l42 = needRd[1];
  always @(*) begin
    if(when_Dispatcher_l42) begin
      freelistRdShuffle_1 = _zz_freelistRdShuffle_1;
    end else begin
      freelistRdShuffle_1 = 6'h00;
    end
  end

  always @(*) begin
    csrReq[0] = (((io_input_availMask[0] && (io_input_dispatchInfo_0_fuType == FUType_csr)) && (! io_aluHasCSRInst_0)) && io_alu0IQ_ready);
    csrReq[1] = (((io_input_availMask[1] && (io_input_dispatchInfo_1_fuType == FUType_csr)) && (! io_aluHasCSRInst_0)) && io_alu0IQ_ready);
  end

  always @(*) begin
    counterReq[0] = (((io_input_availMask[0] && (io_input_dispatchInfo_0_fuType == FUType_counter)) && (! io_aluHasCSRInst_1)) && io_alu1IQ_ready);
    counterReq[1] = (((io_input_availMask[1] && (io_input_dispatchInfo_1_fuType == FUType_counter)) && (! io_aluHasCSRInst_1)) && io_alu1IQ_ready);
  end

  always @(*) begin
    alu0Req[0] = ((io_input_availMask[0] && (io_input_dispatchInfo_0_fuType == FUType_alu)) && io_alu0IQ_ready);
    alu0Req[1] = ((io_input_availMask[1] && (io_input_dispatchInfo_1_fuType == FUType_alu)) && io_alu0IQ_ready);
  end

  always @(*) begin
    alu1Req[0] = ((io_input_availMask[0] && (io_input_dispatchInfo_0_fuType == FUType_alu)) && io_alu1IQ_ready);
    alu1Req[1] = ((io_input_availMask[1] && (io_input_dispatchInfo_1_fuType == FUType_alu)) && io_alu1IQ_ready);
  end

  always @(*) begin
    muluReq[0] = ((io_input_availMask[0] && (io_input_dispatchInfo_0_fuType == FUType_mulu)) && io_muluIQ_ready);
    muluReq[1] = ((io_input_availMask[1] && (io_input_dispatchInfo_1_fuType == FUType_mulu)) && io_muluIQ_ready);
  end

  always @(*) begin
    divuReq[0] = ((io_input_availMask[0] && (io_input_dispatchInfo_0_fuType == FUType_divu)) && io_divuIQ_ready);
    divuReq[1] = ((io_input_availMask[1] && (io_input_dispatchInfo_1_fuType == FUType_divu)) && io_divuIQ_ready);
  end

  always @(*) begin
    lsuReq[0] = ((io_input_availMask[0] && (io_input_dispatchInfo_0_fuType == FUType_lsu)) && io_lsuIQ_ready);
    lsuReq[1] = ((io_input_availMask[1] && (io_input_dispatchInfo_1_fuType == FUType_lsu)) && io_lsuIQ_ready);
  end

  assign _zz_alu0Sel = (csrReq | alu0Req);
  assign alu0Sel = (_zz_alu0Sel & (~ _zz_alu0Sel_1));
  assign _zz_alu1Sel = ((counterReq | alu1Req) & (~ alu0Sel));
  assign alu1Sel = (_zz_alu1Sel & (~ _zz_alu1Sel_1));
  assign muluReq_ohFirst_input = muluReq;
  assign muluReq_ohFirst_masked = (muluReq_ohFirst_input & (~ _zz_muluReq_ohFirst_masked));
  assign muluSel = muluReq_ohFirst_masked;
  assign divuReq_ohFirst_input = divuReq;
  assign divuReq_ohFirst_masked = (divuReq_ohFirst_input & (~ _zz_divuReq_ohFirst_masked));
  assign divuSel = divuReq_ohFirst_masked;
  assign lsuReq_ohFirst_input = lsuReq;
  assign lsuReq_ohFirst_masked = (lsuReq_ohFirst_input & (~ _zz_lsuReq_ohFirst_masked));
  assign lsuSel = lsuReq_ohFirst_masked;
  assign iqAvail = ((((alu0Sel | alu1Sel) | muluSel) | divuSel) | lsuSel);
  assign resAvail = ((freelistAvail & io_rob_availMask) & iqAvail);
  always @(*) begin
    dispatchMask[0] = ((&resAvail[0 : 0]) && io_input_availMask[0]);
    dispatchMask[1] = ((&resAvail[1 : 0]) && io_input_availMask[1]);
  end

  assign io_input_allowMask = dispatchMask;
  assign io_rob_allowMask = dispatchMask;
  assign io_freelist_disPatchNum = _zz_io_freelist_disPatchNum;
  assign actualSrc_0_0 = io_sratReadSrc_0_0_prd;
  assign actualSrcReady_0_0 = (1'b0 ? 1'b0 : io_sratReadSrc_0_0_valid);
  assign actualSrc_0_1 = io_sratReadSrc_0_1_prd;
  assign actualSrcReady_0_1 = (1'b0 ? 1'b0 : io_sratReadSrc_0_1_valid);
  assign actualRd_0 = freelistRdShuffle_0;
  assign actualpRd_0 = io_sratReadPPRD_0_prd;
  always @(*) begin
    _zz_actualSrcReady_1_0[0] = 1'b1;
    _zz_actualSrcReady_1_0[1] = (io_input_dispatchInfo_0_ard == io_input_dispatchInfo_1_asrc_0);
  end

  assign _zz_actualSrc_1_0 = _zz_actualSrcReady_1_0;
  always @(*) begin
    _zz_actualSrc_1_0_1[0] = _zz_actualSrc_1_0[1];
    _zz_actualSrc_1_0_1[1] = _zz_actualSrc_1_0[0];
  end

  assign _zz_actualSrc_1_0_2 = (_zz_actualSrc_1_0_1 & (~ _zz__zz_actualSrc_1_0_2));
  always @(*) begin
    _zz_actualSrc_1_0_3[0] = _zz_actualSrc_1_0_2[1];
    _zz_actualSrc_1_0_3[1] = _zz_actualSrc_1_0_2[0];
  end

  assign actualSrc_1_0 = (_zz_actualSrc_1_0_3[0] ? io_sratReadSrc_1_0_prd : actualRd_0);
  assign actualSrcReady_1_0 = ((|_zz_actualSrcReady_1_0[1 : 1]) ? 1'b0 : io_sratReadSrc_1_0_valid);
  always @(*) begin
    _zz_actualSrcReady_1_1[0] = 1'b1;
    _zz_actualSrcReady_1_1[1] = (io_input_dispatchInfo_0_ard == io_input_dispatchInfo_1_asrc_1);
  end

  assign _zz_actualSrc_1_1 = _zz_actualSrcReady_1_1;
  always @(*) begin
    _zz_actualSrc_1_1_1[0] = _zz_actualSrc_1_1[1];
    _zz_actualSrc_1_1_1[1] = _zz_actualSrc_1_1[0];
  end

  assign _zz_actualSrc_1_1_2 = (_zz_actualSrc_1_1_1 & (~ _zz__zz_actualSrc_1_1_2));
  always @(*) begin
    _zz_actualSrc_1_1_3[0] = _zz_actualSrc_1_1_2[1];
    _zz_actualSrc_1_1_3[1] = _zz_actualSrc_1_1_2[0];
  end

  assign actualSrc_1_1 = (_zz_actualSrc_1_1_3[0] ? io_sratReadSrc_1_1_prd : actualRd_0);
  assign actualSrcReady_1_1 = ((|_zz_actualSrcReady_1_1[1 : 1]) ? 1'b0 : io_sratReadSrc_1_1_valid);
  assign actualRd_1 = freelistRdShuffle_1;
  always @(*) begin
    _zz_actualpRd_1[0] = 1'b1;
    _zz_actualpRd_1[1] = (io_input_dispatchInfo_0_ard == io_input_dispatchInfo_1_ard);
  end

  assign _zz_actualpRd_1_1 = _zz_actualpRd_1;
  always @(*) begin
    _zz_actualpRd_1_2[0] = _zz_actualpRd_1_1[1];
    _zz_actualpRd_1_2[1] = _zz_actualpRd_1_1[0];
  end

  assign _zz_actualpRd_1_3 = (_zz_actualpRd_1_2 & (~ _zz__zz_actualpRd_1_3));
  always @(*) begin
    _zz_actualpRd_1_4[0] = _zz_actualpRd_1_3[1];
    _zz_actualpRd_1_4[1] = _zz_actualpRd_1_3[0];
  end

  assign actualpRd_1 = (_zz_actualpRd_1_4[0] ? io_sratReadPPRD_1_prd : actualRd_0);
  assign alu0Candidate_0_robIdx = io_rob_robIdx_0;
  assign alu1Candidate_0_robIdx = io_rob_robIdx_0;
  assign muluCandidate_0_robIdx = io_rob_robIdx_0;
  assign divuCandidate_0_robIdx = io_rob_robIdx_0;
  assign lsuCandidate_0_robIdx = io_rob_robIdx_0;
  assign alu0Candidate_0_branchInfo_predictPC = decoder_0_io_branchInfo_predictPC;
  assign alu0Candidate_0_branchInfo_predictResult = decoder_0_io_branchInfo_predictResult;
  assign alu1Candidate_0_branchInfo_predictPC = decoder_0_io_branchInfo_predictPC;
  assign alu1Candidate_0_branchInfo_predictResult = decoder_0_io_branchInfo_predictResult;
  assign muluCandidate_0_branchResult_targetPC = decoder_0_io_branchResult_targetPC;
  assign muluCandidate_0_branchResult_branchResult = decoder_0_io_branchResult_branchResult;
  assign muluCandidate_0_branchResult_predictFail = decoder_0_io_branchResult_predictFail;
  assign divuCandidate_0_branchResult_targetPC = decoder_0_io_branchResult_targetPC;
  assign divuCandidate_0_branchResult_branchResult = decoder_0_io_branchResult_branchResult;
  assign divuCandidate_0_branchResult_predictFail = decoder_0_io_branchResult_predictFail;
  assign lsuCandidate_0_branchResult_targetPC = decoder_0_io_branchResult_targetPC;
  assign lsuCandidate_0_branchResult_branchResult = decoder_0_io_branchResult_branchResult;
  assign lsuCandidate_0_branchResult_predictFail = decoder_0_io_branchResult_predictFail;
  assign alu0Candidate_0_exceptionInfo_exception = decoder_0_io_exceptionInfo_exception;
  assign alu0Candidate_0_exceptionInfo_eCode = decoder_0_io_exceptionInfo_eCode;
  assign alu0Candidate_0_exceptionInfo_eSubCode = decoder_0_io_exceptionInfo_eSubCode;
  assign alu1Candidate_0_exceptionInfo_exception = decoder_0_io_exceptionInfo_exception;
  assign alu1Candidate_0_exceptionInfo_eCode = decoder_0_io_exceptionInfo_eCode;
  assign alu1Candidate_0_exceptionInfo_eSubCode = decoder_0_io_exceptionInfo_eSubCode;
  assign muluCandidate_0_exceptionInfo_exception = decoder_0_io_exceptionInfo_exception;
  assign muluCandidate_0_exceptionInfo_eCode = decoder_0_io_exceptionInfo_eCode;
  assign muluCandidate_0_exceptionInfo_eSubCode = decoder_0_io_exceptionInfo_eSubCode;
  assign divuCandidate_0_exceptionInfo_exception = decoder_0_io_exceptionInfo_exception;
  assign divuCandidate_0_exceptionInfo_eCode = decoder_0_io_exceptionInfo_eCode;
  assign divuCandidate_0_exceptionInfo_eSubCode = decoder_0_io_exceptionInfo_eSubCode;
  assign lsuCandidate_0_exceptionInfo_exception = decoder_0_io_exceptionInfo_exception;
  assign lsuCandidate_0_exceptionInfo_eCode = decoder_0_io_exceptionInfo_eCode;
  assign lsuCandidate_0_exceptionInfo_eSubCode = decoder_0_io_exceptionInfo_eSubCode;
  assign alu0Candidate_0_pc = decoder_0_io_pc;
  assign alu1Candidate_0_pc = decoder_0_io_pc;
  assign muluCandidate_0_pc = decoder_0_io_pc;
  assign divuCandidate_0_pc = decoder_0_io_pc;
  assign lsuCandidate_0_pc = decoder_0_io_pc;
  assign alu0Candidate_0_prd = actualRd_0;
  assign alu1Candidate_0_prd = actualRd_0;
  assign muluCandidate_0_prd = actualRd_0;
  assign divuCandidate_0_prd = actualRd_0;
  assign lsuCandidate_0_prd = actualRd_0;
  assign alu0Candidate_0_psrc_0 = actualSrc_0_0;
  assign alu1Candidate_0_psrc_0 = actualSrc_0_0;
  assign muluCandidate_0_psrc_0 = actualSrc_0_0;
  assign divuCandidate_0_psrc_0 = actualSrc_0_0;
  assign lsuCandidate_0_psrc_0 = actualSrc_0_0;
  assign alu0Candidate_0_srcReady_0 = actualSrcReady_0_0;
  assign alu1Candidate_0_srcReady_0 = actualSrcReady_0_0;
  assign muluCandidate_0_srcReady_0 = actualSrcReady_0_0;
  assign divuCandidate_0_srcReady_0 = actualSrcReady_0_0;
  assign lsuCandidate_0_srcReady_0 = actualSrcReady_0_0;
  assign alu0Candidate_0_psrc_1 = actualSrc_0_1;
  assign alu1Candidate_0_psrc_1 = actualSrc_0_1;
  assign muluCandidate_0_psrc_1 = actualSrc_0_1;
  assign divuCandidate_0_psrc_1 = actualSrc_0_1;
  assign lsuCandidate_0_psrc_1 = actualSrc_0_1;
  assign alu0Candidate_0_srcReady_1 = actualSrcReady_0_1;
  assign alu1Candidate_0_srcReady_1 = actualSrcReady_0_1;
  assign muluCandidate_0_srcReady_1 = actualSrcReady_0_1;
  assign divuCandidate_0_srcReady_1 = actualSrcReady_0_1;
  assign lsuCandidate_0_srcReady_1 = actualSrcReady_0_1;
  assign alu0Candidate_0_imm = decoder_0_io_imm;
  assign alu1Candidate_0_imm = decoder_0_io_imm;
  assign muluCandidate_0_imm = decoder_0_io_imm;
  assign divuCandidate_0_imm = decoder_0_io_imm;
  assign lsuCandidate_0_imm = decoder_0_io_imm;
  assign alu0Candidate_0_uop_aluOp = decoder_0_io_uopALU0_aluOp;
  assign alu0Candidate_0_uop_bruOp = decoder_0_io_uopALU0_bruOp;
  assign alu0Candidate_0_uop_cruOp = decoder_0_io_uopALU0_cruOp;
  assign alu1Candidate_0_uop_aluOp = decoder_0_io_uopALU1_aluOp;
  assign alu1Candidate_0_uop_bruOp = decoder_0_io_uopALU1_bruOp;
  assign muluCandidate_0_uop_muluOp = decoder_0_io_uopMULU_muluOp;
  assign divuCandidate_0_uop_divuOp = decoder_0_io_uopDIVU_divuOp;
  assign lsuCandidate_0_uop_lsuOp = decoder_0_io_uopLSU_lsuOp;
  assign lsuCandidate_0_uop_lsuCoOp = decoder_0_io_uopLSU_lsuCoOp;
  assign alu0Candidate_0_roop_aluROOp = decoder_0_io_roopALU0_aluROOp;
  assign alu1Candidate_0_roop_aluROOp = decoder_0_io_roopALU1_aluROOp;
  assign alu1Candidate_0_roop_cruROOp = decoder_0_io_roopALU1_cruROOp;
  assign lsuCandidate_0_roop_lsuROOp = decoder_0_io_roopLSU_lsuROOp;
  assign io_rob_pc_0 = decoder_0_io_pc;
  assign io_rob_ard_0 = io_input_dispatchInfo_0_ard;
  assign io_rob_prd_0 = actualRd_0;
  assign io_rob_pprd_0 = actualpRd_0;
  assign io_rob_specialOp_0 = decoder_0_io_specialOp;
  assign io_sratWrite_0_ard = io_input_dispatchInfo_0_ard;
  assign io_sratWrite_0_prd = actualRd_0;
  assign io_sratWrite_0_wen = (dispatchMask[0] && needRd[0]);
  assign io_sratReadPPRD_0_ard = io_input_dispatchInfo_0_ard;
  assign io_sratReadSrc_0_0_ard = io_input_dispatchInfo_0_asrc_0;
  assign io_sratReadSrc_0_1_ard = io_input_dispatchInfo_0_asrc_1;
  assign alu0Candidate_1_robIdx = io_rob_robIdx_1;
  assign alu1Candidate_1_robIdx = io_rob_robIdx_1;
  assign muluCandidate_1_robIdx = io_rob_robIdx_1;
  assign divuCandidate_1_robIdx = io_rob_robIdx_1;
  assign lsuCandidate_1_robIdx = io_rob_robIdx_1;
  assign alu0Candidate_1_branchInfo_predictPC = decoder_1_1_io_branchInfo_predictPC;
  assign alu0Candidate_1_branchInfo_predictResult = decoder_1_1_io_branchInfo_predictResult;
  assign alu1Candidate_1_branchInfo_predictPC = decoder_1_1_io_branchInfo_predictPC;
  assign alu1Candidate_1_branchInfo_predictResult = decoder_1_1_io_branchInfo_predictResult;
  assign muluCandidate_1_branchResult_targetPC = decoder_1_1_io_branchResult_targetPC;
  assign muluCandidate_1_branchResult_branchResult = decoder_1_1_io_branchResult_branchResult;
  assign muluCandidate_1_branchResult_predictFail = decoder_1_1_io_branchResult_predictFail;
  assign divuCandidate_1_branchResult_targetPC = decoder_1_1_io_branchResult_targetPC;
  assign divuCandidate_1_branchResult_branchResult = decoder_1_1_io_branchResult_branchResult;
  assign divuCandidate_1_branchResult_predictFail = decoder_1_1_io_branchResult_predictFail;
  assign lsuCandidate_1_branchResult_targetPC = decoder_1_1_io_branchResult_targetPC;
  assign lsuCandidate_1_branchResult_branchResult = decoder_1_1_io_branchResult_branchResult;
  assign lsuCandidate_1_branchResult_predictFail = decoder_1_1_io_branchResult_predictFail;
  assign alu0Candidate_1_exceptionInfo_exception = decoder_1_1_io_exceptionInfo_exception;
  assign alu0Candidate_1_exceptionInfo_eCode = decoder_1_1_io_exceptionInfo_eCode;
  assign alu0Candidate_1_exceptionInfo_eSubCode = decoder_1_1_io_exceptionInfo_eSubCode;
  assign alu1Candidate_1_exceptionInfo_exception = decoder_1_1_io_exceptionInfo_exception;
  assign alu1Candidate_1_exceptionInfo_eCode = decoder_1_1_io_exceptionInfo_eCode;
  assign alu1Candidate_1_exceptionInfo_eSubCode = decoder_1_1_io_exceptionInfo_eSubCode;
  assign muluCandidate_1_exceptionInfo_exception = decoder_1_1_io_exceptionInfo_exception;
  assign muluCandidate_1_exceptionInfo_eCode = decoder_1_1_io_exceptionInfo_eCode;
  assign muluCandidate_1_exceptionInfo_eSubCode = decoder_1_1_io_exceptionInfo_eSubCode;
  assign divuCandidate_1_exceptionInfo_exception = decoder_1_1_io_exceptionInfo_exception;
  assign divuCandidate_1_exceptionInfo_eCode = decoder_1_1_io_exceptionInfo_eCode;
  assign divuCandidate_1_exceptionInfo_eSubCode = decoder_1_1_io_exceptionInfo_eSubCode;
  assign lsuCandidate_1_exceptionInfo_exception = decoder_1_1_io_exceptionInfo_exception;
  assign lsuCandidate_1_exceptionInfo_eCode = decoder_1_1_io_exceptionInfo_eCode;
  assign lsuCandidate_1_exceptionInfo_eSubCode = decoder_1_1_io_exceptionInfo_eSubCode;
  assign alu0Candidate_1_pc = decoder_1_1_io_pc;
  assign alu1Candidate_1_pc = decoder_1_1_io_pc;
  assign muluCandidate_1_pc = decoder_1_1_io_pc;
  assign divuCandidate_1_pc = decoder_1_1_io_pc;
  assign lsuCandidate_1_pc = decoder_1_1_io_pc;
  assign alu0Candidate_1_prd = actualRd_1;
  assign alu1Candidate_1_prd = actualRd_1;
  assign muluCandidate_1_prd = actualRd_1;
  assign divuCandidate_1_prd = actualRd_1;
  assign lsuCandidate_1_prd = actualRd_1;
  assign alu0Candidate_1_psrc_0 = actualSrc_1_0;
  assign alu1Candidate_1_psrc_0 = actualSrc_1_0;
  assign muluCandidate_1_psrc_0 = actualSrc_1_0;
  assign divuCandidate_1_psrc_0 = actualSrc_1_0;
  assign lsuCandidate_1_psrc_0 = actualSrc_1_0;
  assign alu0Candidate_1_srcReady_0 = actualSrcReady_1_0;
  assign alu1Candidate_1_srcReady_0 = actualSrcReady_1_0;
  assign muluCandidate_1_srcReady_0 = actualSrcReady_1_0;
  assign divuCandidate_1_srcReady_0 = actualSrcReady_1_0;
  assign lsuCandidate_1_srcReady_0 = actualSrcReady_1_0;
  assign alu0Candidate_1_psrc_1 = actualSrc_1_1;
  assign alu1Candidate_1_psrc_1 = actualSrc_1_1;
  assign muluCandidate_1_psrc_1 = actualSrc_1_1;
  assign divuCandidate_1_psrc_1 = actualSrc_1_1;
  assign lsuCandidate_1_psrc_1 = actualSrc_1_1;
  assign alu0Candidate_1_srcReady_1 = actualSrcReady_1_1;
  assign alu1Candidate_1_srcReady_1 = actualSrcReady_1_1;
  assign muluCandidate_1_srcReady_1 = actualSrcReady_1_1;
  assign divuCandidate_1_srcReady_1 = actualSrcReady_1_1;
  assign lsuCandidate_1_srcReady_1 = actualSrcReady_1_1;
  assign alu0Candidate_1_imm = decoder_1_1_io_imm;
  assign alu1Candidate_1_imm = decoder_1_1_io_imm;
  assign muluCandidate_1_imm = decoder_1_1_io_imm;
  assign divuCandidate_1_imm = decoder_1_1_io_imm;
  assign lsuCandidate_1_imm = decoder_1_1_io_imm;
  assign alu0Candidate_1_uop_aluOp = decoder_1_1_io_uopALU0_aluOp;
  assign alu0Candidate_1_uop_bruOp = decoder_1_1_io_uopALU0_bruOp;
  assign alu0Candidate_1_uop_cruOp = decoder_1_1_io_uopALU0_cruOp;
  assign alu1Candidate_1_uop_aluOp = decoder_1_1_io_uopALU1_aluOp;
  assign alu1Candidate_1_uop_bruOp = decoder_1_1_io_uopALU1_bruOp;
  assign muluCandidate_1_uop_muluOp = decoder_1_1_io_uopMULU_muluOp;
  assign divuCandidate_1_uop_divuOp = decoder_1_1_io_uopDIVU_divuOp;
  assign lsuCandidate_1_uop_lsuOp = decoder_1_1_io_uopLSU_lsuOp;
  assign lsuCandidate_1_uop_lsuCoOp = decoder_1_1_io_uopLSU_lsuCoOp;
  assign alu0Candidate_1_roop_aluROOp = decoder_1_1_io_roopALU0_aluROOp;
  assign alu1Candidate_1_roop_aluROOp = decoder_1_1_io_roopALU1_aluROOp;
  assign alu1Candidate_1_roop_cruROOp = decoder_1_1_io_roopALU1_cruROOp;
  assign lsuCandidate_1_roop_lsuROOp = decoder_1_1_io_roopLSU_lsuROOp;
  assign io_rob_pc_1 = decoder_1_1_io_pc;
  assign io_rob_ard_1 = io_input_dispatchInfo_1_ard;
  assign io_rob_prd_1 = actualRd_1;
  assign io_rob_pprd_1 = actualpRd_1;
  assign io_rob_specialOp_1 = decoder_1_1_io_specialOp;
  assign io_sratWrite_1_ard = io_input_dispatchInfo_1_ard;
  assign io_sratWrite_1_prd = actualRd_1;
  assign io_sratWrite_1_wen = (dispatchMask[1] && needRd[1]);
  assign io_sratReadPPRD_1_ard = io_input_dispatchInfo_1_ard;
  assign io_sratReadSrc_1_0_ard = io_input_dispatchInfo_1_asrc_0;
  assign io_sratReadSrc_1_1_ard = io_input_dispatchInfo_1_asrc_1;
  assign io_alu0IQ_valid = (|(alu0Sel & dispatchMask));
  assign _zz_io_alu0IQ_payload_robIdx = alu0Sel[0];
  assign _zz_io_alu0IQ_payload_uop_aluOp = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_uop_aluOp : alu0Candidate_1_uop_aluOp);
  assign _zz_io_alu0IQ_payload_uop_bruOp = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_uop_bruOp : alu0Candidate_1_uop_bruOp);
  assign _zz_io_alu0IQ_payload_uop_cruOp = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_uop_cruOp : alu0Candidate_1_uop_cruOp);
  assign _zz_io_alu0IQ_payload_roop_aluROOp = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_roop_aluROOp : alu0Candidate_1_roop_aluROOp);
  assign io_alu0IQ_payload_robIdx = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_robIdx : alu0Candidate_1_robIdx);
  assign io_alu0IQ_payload_branchInfo_predictPC = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_branchInfo_predictPC : alu0Candidate_1_branchInfo_predictPC);
  assign io_alu0IQ_payload_branchInfo_predictResult = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_branchInfo_predictResult : alu0Candidate_1_branchInfo_predictResult);
  assign io_alu0IQ_payload_exceptionInfo_exception = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_exceptionInfo_exception : alu0Candidate_1_exceptionInfo_exception);
  assign io_alu0IQ_payload_exceptionInfo_eCode = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_exceptionInfo_eCode : alu0Candidate_1_exceptionInfo_eCode);
  assign io_alu0IQ_payload_exceptionInfo_eSubCode = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_exceptionInfo_eSubCode : alu0Candidate_1_exceptionInfo_eSubCode);
  assign io_alu0IQ_payload_pc = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_pc : alu0Candidate_1_pc);
  assign io_alu0IQ_payload_prd = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_prd : alu0Candidate_1_prd);
  assign io_alu0IQ_payload_psrc_0 = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_psrc_0 : alu0Candidate_1_psrc_0);
  assign io_alu0IQ_payload_psrc_1 = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_psrc_1 : alu0Candidate_1_psrc_1);
  assign io_alu0IQ_payload_imm = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_imm : alu0Candidate_1_imm);
  assign io_alu0IQ_payload_uop_aluOp = _zz_io_alu0IQ_payload_uop_aluOp;
  assign io_alu0IQ_payload_uop_bruOp = _zz_io_alu0IQ_payload_uop_bruOp;
  assign io_alu0IQ_payload_uop_cruOp = _zz_io_alu0IQ_payload_uop_cruOp;
  assign io_alu0IQ_payload_roop_aluROOp = _zz_io_alu0IQ_payload_roop_aluROOp;
  assign io_alu0IQ_payload_srcReady_0 = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_srcReady_0 : alu0Candidate_1_srcReady_0);
  assign io_alu0IQ_payload_srcReady_1 = (_zz_io_alu0IQ_payload_robIdx ? alu0Candidate_0_srcReady_1 : alu0Candidate_1_srcReady_1);
  assign io_alu1IQ_valid = (|(alu1Sel & dispatchMask));
  assign _zz_io_alu1IQ_payload_robIdx = alu1Sel[0];
  assign _zz_io_alu1IQ_payload_uop_aluOp = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_uop_aluOp : alu1Candidate_1_uop_aluOp);
  assign _zz_io_alu1IQ_payload_uop_bruOp = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_uop_bruOp : alu1Candidate_1_uop_bruOp);
  assign _zz_io_alu1IQ_payload_roop_aluROOp = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_roop_aluROOp : alu1Candidate_1_roop_aluROOp);
  assign _zz_io_alu1IQ_payload_roop_cruROOp = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_roop_cruROOp : alu1Candidate_1_roop_cruROOp);
  assign io_alu1IQ_payload_robIdx = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_robIdx : alu1Candidate_1_robIdx);
  assign io_alu1IQ_payload_branchInfo_predictPC = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_branchInfo_predictPC : alu1Candidate_1_branchInfo_predictPC);
  assign io_alu1IQ_payload_branchInfo_predictResult = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_branchInfo_predictResult : alu1Candidate_1_branchInfo_predictResult);
  assign io_alu1IQ_payload_exceptionInfo_exception = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_exceptionInfo_exception : alu1Candidate_1_exceptionInfo_exception);
  assign io_alu1IQ_payload_exceptionInfo_eCode = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_exceptionInfo_eCode : alu1Candidate_1_exceptionInfo_eCode);
  assign io_alu1IQ_payload_exceptionInfo_eSubCode = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_exceptionInfo_eSubCode : alu1Candidate_1_exceptionInfo_eSubCode);
  assign io_alu1IQ_payload_pc = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_pc : alu1Candidate_1_pc);
  assign io_alu1IQ_payload_prd = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_prd : alu1Candidate_1_prd);
  assign io_alu1IQ_payload_psrc_0 = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_psrc_0 : alu1Candidate_1_psrc_0);
  assign io_alu1IQ_payload_psrc_1 = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_psrc_1 : alu1Candidate_1_psrc_1);
  assign io_alu1IQ_payload_imm = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_imm : alu1Candidate_1_imm);
  assign io_alu1IQ_payload_uop_aluOp = _zz_io_alu1IQ_payload_uop_aluOp;
  assign io_alu1IQ_payload_uop_bruOp = _zz_io_alu1IQ_payload_uop_bruOp;
  assign io_alu1IQ_payload_roop_aluROOp = _zz_io_alu1IQ_payload_roop_aluROOp;
  assign io_alu1IQ_payload_roop_cruROOp = _zz_io_alu1IQ_payload_roop_cruROOp;
  assign io_alu1IQ_payload_srcReady_0 = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_srcReady_0 : alu1Candidate_1_srcReady_0);
  assign io_alu1IQ_payload_srcReady_1 = (_zz_io_alu1IQ_payload_robIdx ? alu1Candidate_0_srcReady_1 : alu1Candidate_1_srcReady_1);
  assign io_muluIQ_valid = (|(muluSel & dispatchMask));
  assign _zz_io_muluIQ_payload_robIdx = muluSel[0];
  assign _zz_io_muluIQ_payload_uop_muluOp = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_uop_muluOp : muluCandidate_1_uop_muluOp);
  assign io_muluIQ_payload_robIdx = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_robIdx : muluCandidate_1_robIdx);
  assign io_muluIQ_payload_branchResult_targetPC = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_branchResult_targetPC : muluCandidate_1_branchResult_targetPC);
  assign io_muluIQ_payload_branchResult_branchResult = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_branchResult_branchResult : muluCandidate_1_branchResult_branchResult);
  assign io_muluIQ_payload_branchResult_predictFail = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_branchResult_predictFail : muluCandidate_1_branchResult_predictFail);
  assign io_muluIQ_payload_exceptionInfo_exception = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_exceptionInfo_exception : muluCandidate_1_exceptionInfo_exception);
  assign io_muluIQ_payload_exceptionInfo_eCode = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_exceptionInfo_eCode : muluCandidate_1_exceptionInfo_eCode);
  assign io_muluIQ_payload_exceptionInfo_eSubCode = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_exceptionInfo_eSubCode : muluCandidate_1_exceptionInfo_eSubCode);
  assign io_muluIQ_payload_pc = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_pc : muluCandidate_1_pc);
  assign io_muluIQ_payload_prd = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_prd : muluCandidate_1_prd);
  assign io_muluIQ_payload_psrc_0 = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_psrc_0 : muluCandidate_1_psrc_0);
  assign io_muluIQ_payload_psrc_1 = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_psrc_1 : muluCandidate_1_psrc_1);
  assign io_muluIQ_payload_imm = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_imm : muluCandidate_1_imm);
  assign io_muluIQ_payload_uop_muluOp = _zz_io_muluIQ_payload_uop_muluOp;
  assign io_muluIQ_payload_srcReady_0 = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_srcReady_0 : muluCandidate_1_srcReady_0);
  assign io_muluIQ_payload_srcReady_1 = (_zz_io_muluIQ_payload_robIdx ? muluCandidate_0_srcReady_1 : muluCandidate_1_srcReady_1);
  assign io_divuIQ_valid = (|(divuSel & dispatchMask));
  assign _zz_io_divuIQ_payload_robIdx = divuSel[0];
  assign _zz_io_divuIQ_payload_uop_divuOp = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_uop_divuOp : divuCandidate_1_uop_divuOp);
  assign io_divuIQ_payload_robIdx = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_robIdx : divuCandidate_1_robIdx);
  assign io_divuIQ_payload_branchResult_targetPC = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_branchResult_targetPC : divuCandidate_1_branchResult_targetPC);
  assign io_divuIQ_payload_branchResult_branchResult = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_branchResult_branchResult : divuCandidate_1_branchResult_branchResult);
  assign io_divuIQ_payload_branchResult_predictFail = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_branchResult_predictFail : divuCandidate_1_branchResult_predictFail);
  assign io_divuIQ_payload_exceptionInfo_exception = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_exceptionInfo_exception : divuCandidate_1_exceptionInfo_exception);
  assign io_divuIQ_payload_exceptionInfo_eCode = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_exceptionInfo_eCode : divuCandidate_1_exceptionInfo_eCode);
  assign io_divuIQ_payload_exceptionInfo_eSubCode = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_exceptionInfo_eSubCode : divuCandidate_1_exceptionInfo_eSubCode);
  assign io_divuIQ_payload_pc = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_pc : divuCandidate_1_pc);
  assign io_divuIQ_payload_prd = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_prd : divuCandidate_1_prd);
  assign io_divuIQ_payload_psrc_0 = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_psrc_0 : divuCandidate_1_psrc_0);
  assign io_divuIQ_payload_psrc_1 = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_psrc_1 : divuCandidate_1_psrc_1);
  assign io_divuIQ_payload_imm = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_imm : divuCandidate_1_imm);
  assign io_divuIQ_payload_uop_divuOp = _zz_io_divuIQ_payload_uop_divuOp;
  assign io_divuIQ_payload_srcReady_0 = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_srcReady_0 : divuCandidate_1_srcReady_0);
  assign io_divuIQ_payload_srcReady_1 = (_zz_io_divuIQ_payload_robIdx ? divuCandidate_0_srcReady_1 : divuCandidate_1_srcReady_1);
  assign io_lsuIQ_valid = (|(lsuSel & dispatchMask));
  assign _zz_io_lsuIQ_payload_robIdx = lsuSel[0];
  assign _zz_io_lsuIQ_payload_uop_lsuOp = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_uop_lsuOp : lsuCandidate_1_uop_lsuOp);
  assign _zz_io_lsuIQ_payload_roop_lsuROOp = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_roop_lsuROOp : lsuCandidate_1_roop_lsuROOp);
  assign io_lsuIQ_payload_robIdx = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_robIdx : lsuCandidate_1_robIdx);
  assign io_lsuIQ_payload_branchResult_targetPC = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_branchResult_targetPC : lsuCandidate_1_branchResult_targetPC);
  assign io_lsuIQ_payload_branchResult_branchResult = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_branchResult_branchResult : lsuCandidate_1_branchResult_branchResult);
  assign io_lsuIQ_payload_branchResult_predictFail = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_branchResult_predictFail : lsuCandidate_1_branchResult_predictFail);
  assign io_lsuIQ_payload_exceptionInfo_exception = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_exceptionInfo_exception : lsuCandidate_1_exceptionInfo_exception);
  assign io_lsuIQ_payload_exceptionInfo_eCode = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_exceptionInfo_eCode : lsuCandidate_1_exceptionInfo_eCode);
  assign io_lsuIQ_payload_exceptionInfo_eSubCode = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_exceptionInfo_eSubCode : lsuCandidate_1_exceptionInfo_eSubCode);
  assign io_lsuIQ_payload_pc = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_pc : lsuCandidate_1_pc);
  assign io_lsuIQ_payload_prd = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_prd : lsuCandidate_1_prd);
  assign io_lsuIQ_payload_psrc_0 = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_psrc_0 : lsuCandidate_1_psrc_0);
  assign io_lsuIQ_payload_psrc_1 = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_psrc_1 : lsuCandidate_1_psrc_1);
  assign io_lsuIQ_payload_imm = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_imm : lsuCandidate_1_imm);
  assign io_lsuIQ_payload_uop_lsuOp = _zz_io_lsuIQ_payload_uop_lsuOp;
  assign io_lsuIQ_payload_uop_lsuCoOp = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_uop_lsuCoOp : lsuCandidate_1_uop_lsuCoOp);
  assign io_lsuIQ_payload_roop_lsuROOp = _zz_io_lsuIQ_payload_roop_lsuROOp;
  assign io_lsuIQ_payload_srcReady_0 = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_srcReady_0 : lsuCandidate_1_srcReady_0);
  assign io_lsuIQ_payload_srcReady_1 = (_zz_io_lsuIQ_payload_robIdx ? lsuCandidate_0_srcReady_1 : lsuCandidate_1_srcReady_1);

endmodule

module InstrQueue (
  output wire [1:0]    io_in_allowMask,
  input  wire [1:0]    io_in_availMask,
  input  wire [31:0]   io_in_info_0_inst,
  input  wire [31:0]   io_in_info_0_branchInfo_predictPC,
  input  wire          io_in_info_0_branchInfo_predictResult,
  input  wire          io_in_info_0_exceptionInfo_exception,
  input  wire [5:0]    io_in_info_0_exceptionInfo_eCode,
  input  wire [0:0]    io_in_info_0_exceptionInfo_eSubCode,
  input  wire [31:0]   io_in_info_0_pc,
  input  wire [31:0]   io_in_info_1_inst,
  input  wire [31:0]   io_in_info_1_branchInfo_predictPC,
  input  wire          io_in_info_1_branchInfo_predictResult,
  input  wire          io_in_info_1_exceptionInfo_exception,
  input  wire [5:0]    io_in_info_1_exceptionInfo_eCode,
  input  wire [0:0]    io_in_info_1_exceptionInfo_eSubCode,
  input  wire [31:0]   io_in_info_1_pc,
  input  wire [1:0]    io_out_allowMask,
  output reg  [1:0]    io_out_availMask,
  output wire [31:0]   io_out_info_0_inst,
  output wire [31:0]   io_out_info_0_branchInfo_predictPC,
  output wire          io_out_info_0_branchInfo_predictResult,
  output wire          io_out_info_0_exceptionInfo_exception,
  output wire [5:0]    io_out_info_0_exceptionInfo_eCode,
  output wire [0:0]    io_out_info_0_exceptionInfo_eSubCode,
  output wire [31:0]   io_out_info_0_pc,
  output wire [31:0]   io_out_info_1_inst,
  output wire [31:0]   io_out_info_1_branchInfo_predictPC,
  output wire          io_out_info_1_branchInfo_predictResult,
  output wire          io_out_info_1_exceptionInfo_exception,
  output wire [5:0]    io_out_info_1_exceptionInfo_eCode,
  output wire [0:0]    io_out_info_1_exceptionInfo_eSubCode,
  output wire [31:0]   io_out_info_1_pc,
  output wire [2:0]    io_out_dispatchInfo_0_fuType,
  output wire [4:0]    io_out_dispatchInfo_0_ard,
  output wire [4:0]    io_out_dispatchInfo_0_asrc_0,
  output wire [4:0]    io_out_dispatchInfo_0_asrc_1,
  output wire [2:0]    io_out_dispatchInfo_1_fuType,
  output wire [4:0]    io_out_dispatchInfo_1_ard,
  output wire [4:0]    io_out_dispatchInfo_1_asrc_0,
  output wire [4:0]    io_out_dispatchInfo_1_asrc_1,
  input  wire          aclk,
  input  wire          cpuClockingArea_areaFlushReset_newReset
);
  localparam FUType_alu = 3'd0;
  localparam FUType_csr = 3'd1;
  localparam FUType_counter = 3'd2;
  localparam FUType_lsu = 3'd3;
  localparam FUType_mulu = 3'd4;
  localparam FUType_divu = 3'd5;

  reg        [1:0]    _zz_fetchNum;
  wire       [1:0]    _zz_fetchNum_1;
  reg        [1:0]    _zz_dispatchNum;
  wire       [1:0]    _zz_dispatchNum_1;
  reg                 _zz_allowMask;
  wire       [2:0]    _zz_tail_0;
  reg                 _zz_allowMask_1;
  wire       [2:0]    _zz_tail_1;
  reg        [31:0]   _zz__zz_io_out_info_0_inst;
  reg        [31:0]   _zz_io_out_info_0_branchInfo_predictPC;
  reg                 _zz_io_out_info_0_branchInfo_predictResult;
  reg                 _zz_io_out_info_0_exceptionInfo_exception;
  reg        [5:0]    _zz_io_out_info_0_exceptionInfo_eCode;
  reg        [0:0]    _zz_io_out_info_0_exceptionInfo_eSubCode;
  reg        [31:0]   _zz_io_out_info_0_pc;
  wire       [0:0]    _zz__zz_io_out_dispatchInfo_0_ard;
  wire       [4:0]    _zz_when_InstrQueue_l119_2;
  wire       [0:0]    _zz_when_InstrQueue_l119_3;
  reg                 _zz_io_out_availMask;
  wire       [2:0]    _zz_head_0;
  reg        [31:0]   _zz__zz_io_out_info_1_inst;
  reg        [31:0]   _zz_io_out_info_1_branchInfo_predictPC;
  reg                 _zz_io_out_info_1_branchInfo_predictResult;
  reg                 _zz_io_out_info_1_exceptionInfo_exception;
  reg        [5:0]    _zz_io_out_info_1_exceptionInfo_eCode;
  reg        [0:0]    _zz_io_out_info_1_exceptionInfo_eSubCode;
  reg        [31:0]   _zz_io_out_info_1_pc;
  wire       [0:0]    _zz__zz_io_out_dispatchInfo_1_ard;
  wire       [4:0]    _zz_when_InstrQueue_l119_1_1;
  wire       [0:0]    _zz_when_InstrQueue_l119_1_2;
  reg                 _zz_io_out_availMask_1;
  wire       [2:0]    _zz_head_1;
  reg        [31:0]   queue_0_inst;
  reg        [31:0]   queue_0_branchInfo_predictPC;
  reg                 queue_0_branchInfo_predictResult;
  reg                 queue_0_exceptionInfo_exception;
  reg        [5:0]    queue_0_exceptionInfo_eCode;
  reg        [0:0]    queue_0_exceptionInfo_eSubCode;
  reg        [31:0]   queue_0_pc;
  reg        [31:0]   queue_1_inst;
  reg        [31:0]   queue_1_branchInfo_predictPC;
  reg                 queue_1_branchInfo_predictResult;
  reg                 queue_1_exceptionInfo_exception;
  reg        [5:0]    queue_1_exceptionInfo_eCode;
  reg        [0:0]    queue_1_exceptionInfo_eSubCode;
  reg        [31:0]   queue_1_pc;
  reg        [31:0]   queue_2_inst;
  reg        [31:0]   queue_2_branchInfo_predictPC;
  reg                 queue_2_branchInfo_predictResult;
  reg                 queue_2_exceptionInfo_exception;
  reg        [5:0]    queue_2_exceptionInfo_eCode;
  reg        [0:0]    queue_2_exceptionInfo_eSubCode;
  reg        [31:0]   queue_2_pc;
  reg        [31:0]   queue_3_inst;
  reg        [31:0]   queue_3_branchInfo_predictPC;
  reg                 queue_3_branchInfo_predictResult;
  reg                 queue_3_exceptionInfo_exception;
  reg        [5:0]    queue_3_exceptionInfo_eCode;
  reg        [0:0]    queue_3_exceptionInfo_eSubCode;
  reg        [31:0]   queue_3_pc;
  reg        [31:0]   queue_4_inst;
  reg        [31:0]   queue_4_branchInfo_predictPC;
  reg                 queue_4_branchInfo_predictResult;
  reg                 queue_4_exceptionInfo_exception;
  reg        [5:0]    queue_4_exceptionInfo_eCode;
  reg        [0:0]    queue_4_exceptionInfo_eSubCode;
  reg        [31:0]   queue_4_pc;
  reg        [31:0]   queue_5_inst;
  reg        [31:0]   queue_5_branchInfo_predictPC;
  reg                 queue_5_branchInfo_predictResult;
  reg                 queue_5_exceptionInfo_exception;
  reg        [5:0]    queue_5_exceptionInfo_eCode;
  reg        [0:0]    queue_5_exceptionInfo_eSubCode;
  reg        [31:0]   queue_5_pc;
  reg        [31:0]   queue_6_inst;
  reg        [31:0]   queue_6_branchInfo_predictPC;
  reg                 queue_6_branchInfo_predictResult;
  reg                 queue_6_exceptionInfo_exception;
  reg        [5:0]    queue_6_exceptionInfo_eCode;
  reg        [0:0]    queue_6_exceptionInfo_eSubCode;
  reg        [31:0]   queue_6_pc;
  reg        [31:0]   queue_7_inst;
  reg        [31:0]   queue_7_branchInfo_predictPC;
  reg                 queue_7_branchInfo_predictResult;
  reg                 queue_7_exceptionInfo_exception;
  reg        [5:0]    queue_7_exceptionInfo_eCode;
  reg        [0:0]    queue_7_exceptionInfo_eSubCode;
  reg        [31:0]   queue_7_pc;
  reg                 valid_0;
  reg                 valid_1;
  reg                 valid_2;
  reg                 valid_3;
  reg                 valid_4;
  reg                 valid_5;
  reg                 valid_6;
  reg                 valid_7;
  reg        [2:0]    head_0;
  reg        [2:0]    head_1;
  reg        [2:0]    tail_0;
  reg        [2:0]    tail_1;
  wire       [1:0]    fetchNum;
  wire       [1:0]    dispatchNum;
  reg        [1:0]    allowMask;
  wire                when_InstrQueue_l33;
  wire       [7:0]    _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                when_InstrQueue_l33_1;
  wire       [7:0]    _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire       [31:0]   _zz_io_out_info_0_inst;
  reg        [2:0]    _zz_io_out_dispatchInfo_0_fuType;
  reg        [4:0]    _zz_io_out_dispatchInfo_0_ard;
  reg        [4:0]    _zz_io_out_dispatchInfo_0_asrc_0;
  reg        [4:0]    _zz_io_out_dispatchInfo_0_asrc_1;
  wire       [4:0]    _zz_io_out_dispatchInfo_0_ard_1;
  wire       [4:0]    _zz_when_InstrQueue_l119;
  wire       [4:0]    _zz_io_out_dispatchInfo_0_asrc_1_1;
  wire       [0:0]    _zz_io_out_dispatchInfo_0_ard_2;
  wire                when_InstrQueue_l119;
  wire       [31:0]   _zz_io_out_info_1_inst;
  reg        [2:0]    _zz_io_out_dispatchInfo_1_fuType;
  reg        [4:0]    _zz_io_out_dispatchInfo_1_ard;
  reg        [4:0]    _zz_io_out_dispatchInfo_1_asrc_0;
  reg        [4:0]    _zz_io_out_dispatchInfo_1_asrc_1;
  wire       [4:0]    _zz_io_out_dispatchInfo_1_ard_1;
  wire       [4:0]    _zz_when_InstrQueue_l119_1;
  wire       [4:0]    _zz_io_out_dispatchInfo_1_asrc_1_1;
  wire       [0:0]    _zz_io_out_dispatchInfo_1_ard_2;
  wire                when_InstrQueue_l119_1;
  reg        [1:0]    _zz_valid_0;
  reg        [1:0]    _zz_valid_0_1;
  reg        [1:0]    _zz_valid_1;
  reg        [1:0]    _zz_valid_1_1;
  reg        [1:0]    _zz_valid_2;
  reg        [1:0]    _zz_valid_2_1;
  reg        [1:0]    _zz_valid_3;
  reg        [1:0]    _zz_valid_3_1;
  reg        [1:0]    _zz_valid_4;
  reg        [1:0]    _zz_valid_4_1;
  reg        [1:0]    _zz_valid_5;
  reg        [1:0]    _zz_valid_5_1;
  reg        [1:0]    _zz_valid_6;
  reg        [1:0]    _zz_valid_6_1;
  reg        [1:0]    _zz_valid_7;
  reg        [1:0]    _zz_valid_7_1;
  `ifndef SYNTHESIS
  reg [55:0] io_out_dispatchInfo_0_fuType_string;
  reg [55:0] io_out_dispatchInfo_1_fuType_string;
  reg [55:0] _zz_io_out_dispatchInfo_0_fuType_string;
  reg [55:0] _zz_io_out_dispatchInfo_1_fuType_string;
  `endif


  assign _zz_tail_0 = {1'd0, fetchNum};
  assign _zz_tail_1 = {1'd0, fetchNum};
  assign _zz__zz_io_out_dispatchInfo_0_ard = 1'b1;
  assign _zz_when_InstrQueue_l119_3 = 1'b1;
  assign _zz_when_InstrQueue_l119_2 = {4'd0, _zz_when_InstrQueue_l119_3};
  assign _zz_head_0 = {1'd0, dispatchNum};
  assign _zz__zz_io_out_dispatchInfo_1_ard = 1'b1;
  assign _zz_when_InstrQueue_l119_1_2 = 1'b1;
  assign _zz_when_InstrQueue_l119_1_1 = {4'd0, _zz_when_InstrQueue_l119_1_2};
  assign _zz_head_1 = {1'd0, dispatchNum};
  assign _zz_fetchNum_1 = {io_in_allowMask[1],io_in_allowMask[0]};
  assign _zz_dispatchNum_1 = {io_out_allowMask[1],io_out_allowMask[0]};
  always @(*) begin
    case(_zz_fetchNum_1)
      2'b00 : _zz_fetchNum = 2'b00;
      2'b01 : _zz_fetchNum = 2'b01;
      2'b10 : _zz_fetchNum = 2'b01;
      default : _zz_fetchNum = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_dispatchNum_1)
      2'b00 : _zz_dispatchNum = 2'b00;
      2'b01 : _zz_dispatchNum = 2'b01;
      2'b10 : _zz_dispatchNum = 2'b01;
      default : _zz_dispatchNum = 2'b10;
    endcase
  end

  always @(*) begin
    case(tail_0)
      3'b000 : _zz_allowMask = valid_0;
      3'b001 : _zz_allowMask = valid_1;
      3'b010 : _zz_allowMask = valid_2;
      3'b011 : _zz_allowMask = valid_3;
      3'b100 : _zz_allowMask = valid_4;
      3'b101 : _zz_allowMask = valid_5;
      3'b110 : _zz_allowMask = valid_6;
      default : _zz_allowMask = valid_7;
    endcase
  end

  always @(*) begin
    case(tail_1)
      3'b000 : _zz_allowMask_1 = valid_0;
      3'b001 : _zz_allowMask_1 = valid_1;
      3'b010 : _zz_allowMask_1 = valid_2;
      3'b011 : _zz_allowMask_1 = valid_3;
      3'b100 : _zz_allowMask_1 = valid_4;
      3'b101 : _zz_allowMask_1 = valid_5;
      3'b110 : _zz_allowMask_1 = valid_6;
      default : _zz_allowMask_1 = valid_7;
    endcase
  end

  always @(*) begin
    case(head_0)
      3'b000 : begin
        _zz__zz_io_out_info_0_inst = queue_0_inst;
        _zz_io_out_info_0_branchInfo_predictPC = queue_0_branchInfo_predictPC;
        _zz_io_out_info_0_branchInfo_predictResult = queue_0_branchInfo_predictResult;
        _zz_io_out_info_0_exceptionInfo_exception = queue_0_exceptionInfo_exception;
        _zz_io_out_info_0_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
        _zz_io_out_info_0_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
        _zz_io_out_info_0_pc = queue_0_pc;
        _zz_io_out_availMask = valid_0;
      end
      3'b001 : begin
        _zz__zz_io_out_info_0_inst = queue_1_inst;
        _zz_io_out_info_0_branchInfo_predictPC = queue_1_branchInfo_predictPC;
        _zz_io_out_info_0_branchInfo_predictResult = queue_1_branchInfo_predictResult;
        _zz_io_out_info_0_exceptionInfo_exception = queue_1_exceptionInfo_exception;
        _zz_io_out_info_0_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
        _zz_io_out_info_0_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
        _zz_io_out_info_0_pc = queue_1_pc;
        _zz_io_out_availMask = valid_1;
      end
      3'b010 : begin
        _zz__zz_io_out_info_0_inst = queue_2_inst;
        _zz_io_out_info_0_branchInfo_predictPC = queue_2_branchInfo_predictPC;
        _zz_io_out_info_0_branchInfo_predictResult = queue_2_branchInfo_predictResult;
        _zz_io_out_info_0_exceptionInfo_exception = queue_2_exceptionInfo_exception;
        _zz_io_out_info_0_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
        _zz_io_out_info_0_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
        _zz_io_out_info_0_pc = queue_2_pc;
        _zz_io_out_availMask = valid_2;
      end
      3'b011 : begin
        _zz__zz_io_out_info_0_inst = queue_3_inst;
        _zz_io_out_info_0_branchInfo_predictPC = queue_3_branchInfo_predictPC;
        _zz_io_out_info_0_branchInfo_predictResult = queue_3_branchInfo_predictResult;
        _zz_io_out_info_0_exceptionInfo_exception = queue_3_exceptionInfo_exception;
        _zz_io_out_info_0_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
        _zz_io_out_info_0_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
        _zz_io_out_info_0_pc = queue_3_pc;
        _zz_io_out_availMask = valid_3;
      end
      3'b100 : begin
        _zz__zz_io_out_info_0_inst = queue_4_inst;
        _zz_io_out_info_0_branchInfo_predictPC = queue_4_branchInfo_predictPC;
        _zz_io_out_info_0_branchInfo_predictResult = queue_4_branchInfo_predictResult;
        _zz_io_out_info_0_exceptionInfo_exception = queue_4_exceptionInfo_exception;
        _zz_io_out_info_0_exceptionInfo_eCode = queue_4_exceptionInfo_eCode;
        _zz_io_out_info_0_exceptionInfo_eSubCode = queue_4_exceptionInfo_eSubCode;
        _zz_io_out_info_0_pc = queue_4_pc;
        _zz_io_out_availMask = valid_4;
      end
      3'b101 : begin
        _zz__zz_io_out_info_0_inst = queue_5_inst;
        _zz_io_out_info_0_branchInfo_predictPC = queue_5_branchInfo_predictPC;
        _zz_io_out_info_0_branchInfo_predictResult = queue_5_branchInfo_predictResult;
        _zz_io_out_info_0_exceptionInfo_exception = queue_5_exceptionInfo_exception;
        _zz_io_out_info_0_exceptionInfo_eCode = queue_5_exceptionInfo_eCode;
        _zz_io_out_info_0_exceptionInfo_eSubCode = queue_5_exceptionInfo_eSubCode;
        _zz_io_out_info_0_pc = queue_5_pc;
        _zz_io_out_availMask = valid_5;
      end
      3'b110 : begin
        _zz__zz_io_out_info_0_inst = queue_6_inst;
        _zz_io_out_info_0_branchInfo_predictPC = queue_6_branchInfo_predictPC;
        _zz_io_out_info_0_branchInfo_predictResult = queue_6_branchInfo_predictResult;
        _zz_io_out_info_0_exceptionInfo_exception = queue_6_exceptionInfo_exception;
        _zz_io_out_info_0_exceptionInfo_eCode = queue_6_exceptionInfo_eCode;
        _zz_io_out_info_0_exceptionInfo_eSubCode = queue_6_exceptionInfo_eSubCode;
        _zz_io_out_info_0_pc = queue_6_pc;
        _zz_io_out_availMask = valid_6;
      end
      default : begin
        _zz__zz_io_out_info_0_inst = queue_7_inst;
        _zz_io_out_info_0_branchInfo_predictPC = queue_7_branchInfo_predictPC;
        _zz_io_out_info_0_branchInfo_predictResult = queue_7_branchInfo_predictResult;
        _zz_io_out_info_0_exceptionInfo_exception = queue_7_exceptionInfo_exception;
        _zz_io_out_info_0_exceptionInfo_eCode = queue_7_exceptionInfo_eCode;
        _zz_io_out_info_0_exceptionInfo_eSubCode = queue_7_exceptionInfo_eSubCode;
        _zz_io_out_info_0_pc = queue_7_pc;
        _zz_io_out_availMask = valid_7;
      end
    endcase
  end

  always @(*) begin
    case(head_1)
      3'b000 : begin
        _zz__zz_io_out_info_1_inst = queue_0_inst;
        _zz_io_out_info_1_branchInfo_predictPC = queue_0_branchInfo_predictPC;
        _zz_io_out_info_1_branchInfo_predictResult = queue_0_branchInfo_predictResult;
        _zz_io_out_info_1_exceptionInfo_exception = queue_0_exceptionInfo_exception;
        _zz_io_out_info_1_exceptionInfo_eCode = queue_0_exceptionInfo_eCode;
        _zz_io_out_info_1_exceptionInfo_eSubCode = queue_0_exceptionInfo_eSubCode;
        _zz_io_out_info_1_pc = queue_0_pc;
        _zz_io_out_availMask_1 = valid_0;
      end
      3'b001 : begin
        _zz__zz_io_out_info_1_inst = queue_1_inst;
        _zz_io_out_info_1_branchInfo_predictPC = queue_1_branchInfo_predictPC;
        _zz_io_out_info_1_branchInfo_predictResult = queue_1_branchInfo_predictResult;
        _zz_io_out_info_1_exceptionInfo_exception = queue_1_exceptionInfo_exception;
        _zz_io_out_info_1_exceptionInfo_eCode = queue_1_exceptionInfo_eCode;
        _zz_io_out_info_1_exceptionInfo_eSubCode = queue_1_exceptionInfo_eSubCode;
        _zz_io_out_info_1_pc = queue_1_pc;
        _zz_io_out_availMask_1 = valid_1;
      end
      3'b010 : begin
        _zz__zz_io_out_info_1_inst = queue_2_inst;
        _zz_io_out_info_1_branchInfo_predictPC = queue_2_branchInfo_predictPC;
        _zz_io_out_info_1_branchInfo_predictResult = queue_2_branchInfo_predictResult;
        _zz_io_out_info_1_exceptionInfo_exception = queue_2_exceptionInfo_exception;
        _zz_io_out_info_1_exceptionInfo_eCode = queue_2_exceptionInfo_eCode;
        _zz_io_out_info_1_exceptionInfo_eSubCode = queue_2_exceptionInfo_eSubCode;
        _zz_io_out_info_1_pc = queue_2_pc;
        _zz_io_out_availMask_1 = valid_2;
      end
      3'b011 : begin
        _zz__zz_io_out_info_1_inst = queue_3_inst;
        _zz_io_out_info_1_branchInfo_predictPC = queue_3_branchInfo_predictPC;
        _zz_io_out_info_1_branchInfo_predictResult = queue_3_branchInfo_predictResult;
        _zz_io_out_info_1_exceptionInfo_exception = queue_3_exceptionInfo_exception;
        _zz_io_out_info_1_exceptionInfo_eCode = queue_3_exceptionInfo_eCode;
        _zz_io_out_info_1_exceptionInfo_eSubCode = queue_3_exceptionInfo_eSubCode;
        _zz_io_out_info_1_pc = queue_3_pc;
        _zz_io_out_availMask_1 = valid_3;
      end
      3'b100 : begin
        _zz__zz_io_out_info_1_inst = queue_4_inst;
        _zz_io_out_info_1_branchInfo_predictPC = queue_4_branchInfo_predictPC;
        _zz_io_out_info_1_branchInfo_predictResult = queue_4_branchInfo_predictResult;
        _zz_io_out_info_1_exceptionInfo_exception = queue_4_exceptionInfo_exception;
        _zz_io_out_info_1_exceptionInfo_eCode = queue_4_exceptionInfo_eCode;
        _zz_io_out_info_1_exceptionInfo_eSubCode = queue_4_exceptionInfo_eSubCode;
        _zz_io_out_info_1_pc = queue_4_pc;
        _zz_io_out_availMask_1 = valid_4;
      end
      3'b101 : begin
        _zz__zz_io_out_info_1_inst = queue_5_inst;
        _zz_io_out_info_1_branchInfo_predictPC = queue_5_branchInfo_predictPC;
        _zz_io_out_info_1_branchInfo_predictResult = queue_5_branchInfo_predictResult;
        _zz_io_out_info_1_exceptionInfo_exception = queue_5_exceptionInfo_exception;
        _zz_io_out_info_1_exceptionInfo_eCode = queue_5_exceptionInfo_eCode;
        _zz_io_out_info_1_exceptionInfo_eSubCode = queue_5_exceptionInfo_eSubCode;
        _zz_io_out_info_1_pc = queue_5_pc;
        _zz_io_out_availMask_1 = valid_5;
      end
      3'b110 : begin
        _zz__zz_io_out_info_1_inst = queue_6_inst;
        _zz_io_out_info_1_branchInfo_predictPC = queue_6_branchInfo_predictPC;
        _zz_io_out_info_1_branchInfo_predictResult = queue_6_branchInfo_predictResult;
        _zz_io_out_info_1_exceptionInfo_exception = queue_6_exceptionInfo_exception;
        _zz_io_out_info_1_exceptionInfo_eCode = queue_6_exceptionInfo_eCode;
        _zz_io_out_info_1_exceptionInfo_eSubCode = queue_6_exceptionInfo_eSubCode;
        _zz_io_out_info_1_pc = queue_6_pc;
        _zz_io_out_availMask_1 = valid_6;
      end
      default : begin
        _zz__zz_io_out_info_1_inst = queue_7_inst;
        _zz_io_out_info_1_branchInfo_predictPC = queue_7_branchInfo_predictPC;
        _zz_io_out_info_1_branchInfo_predictResult = queue_7_branchInfo_predictResult;
        _zz_io_out_info_1_exceptionInfo_exception = queue_7_exceptionInfo_exception;
        _zz_io_out_info_1_exceptionInfo_eCode = queue_7_exceptionInfo_eCode;
        _zz_io_out_info_1_exceptionInfo_eSubCode = queue_7_exceptionInfo_eSubCode;
        _zz_io_out_info_1_pc = queue_7_pc;
        _zz_io_out_availMask_1 = valid_7;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_out_dispatchInfo_0_fuType)
      FUType_alu : io_out_dispatchInfo_0_fuType_string = "alu    ";
      FUType_csr : io_out_dispatchInfo_0_fuType_string = "csr    ";
      FUType_counter : io_out_dispatchInfo_0_fuType_string = "counter";
      FUType_lsu : io_out_dispatchInfo_0_fuType_string = "lsu    ";
      FUType_mulu : io_out_dispatchInfo_0_fuType_string = "mulu   ";
      FUType_divu : io_out_dispatchInfo_0_fuType_string = "divu   ";
      default : io_out_dispatchInfo_0_fuType_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_out_dispatchInfo_1_fuType)
      FUType_alu : io_out_dispatchInfo_1_fuType_string = "alu    ";
      FUType_csr : io_out_dispatchInfo_1_fuType_string = "csr    ";
      FUType_counter : io_out_dispatchInfo_1_fuType_string = "counter";
      FUType_lsu : io_out_dispatchInfo_1_fuType_string = "lsu    ";
      FUType_mulu : io_out_dispatchInfo_1_fuType_string = "mulu   ";
      FUType_divu : io_out_dispatchInfo_1_fuType_string = "divu   ";
      default : io_out_dispatchInfo_1_fuType_string = "???????";
    endcase
  end
  always @(*) begin
    case(_zz_io_out_dispatchInfo_0_fuType)
      FUType_alu : _zz_io_out_dispatchInfo_0_fuType_string = "alu    ";
      FUType_csr : _zz_io_out_dispatchInfo_0_fuType_string = "csr    ";
      FUType_counter : _zz_io_out_dispatchInfo_0_fuType_string = "counter";
      FUType_lsu : _zz_io_out_dispatchInfo_0_fuType_string = "lsu    ";
      FUType_mulu : _zz_io_out_dispatchInfo_0_fuType_string = "mulu   ";
      FUType_divu : _zz_io_out_dispatchInfo_0_fuType_string = "divu   ";
      default : _zz_io_out_dispatchInfo_0_fuType_string = "???????";
    endcase
  end
  always @(*) begin
    case(_zz_io_out_dispatchInfo_1_fuType)
      FUType_alu : _zz_io_out_dispatchInfo_1_fuType_string = "alu    ";
      FUType_csr : _zz_io_out_dispatchInfo_1_fuType_string = "csr    ";
      FUType_counter : _zz_io_out_dispatchInfo_1_fuType_string = "counter";
      FUType_lsu : _zz_io_out_dispatchInfo_1_fuType_string = "lsu    ";
      FUType_mulu : _zz_io_out_dispatchInfo_1_fuType_string = "mulu   ";
      FUType_divu : _zz_io_out_dispatchInfo_1_fuType_string = "divu   ";
      default : _zz_io_out_dispatchInfo_1_fuType_string = "???????";
    endcase
  end
  `endif

  assign fetchNum = _zz_fetchNum;
  assign dispatchNum = _zz_dispatchNum;
  assign io_in_allowMask = (allowMask & io_in_availMask);
  always @(*) begin
    allowMask[0] = (! _zz_allowMask);
    allowMask[1] = (! _zz_allowMask_1);
  end

  assign when_InstrQueue_l33 = io_in_allowMask[0];
  assign _zz_1 = ({7'd0,1'b1} <<< tail_0);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = _zz_1[4];
  assign _zz_7 = _zz_1[5];
  assign _zz_8 = _zz_1[6];
  assign _zz_9 = _zz_1[7];
  assign when_InstrQueue_l33_1 = io_in_allowMask[1];
  assign _zz_10 = ({7'd0,1'b1} <<< tail_1);
  assign _zz_11 = _zz_10[0];
  assign _zz_12 = _zz_10[1];
  assign _zz_13 = _zz_10[2];
  assign _zz_14 = _zz_10[3];
  assign _zz_15 = _zz_10[4];
  assign _zz_16 = _zz_10[5];
  assign _zz_17 = _zz_10[6];
  assign _zz_18 = _zz_10[7];
  assign _zz_io_out_info_0_inst = _zz__zz_io_out_info_0_inst;
  assign io_out_info_0_inst = _zz_io_out_info_0_inst;
  assign io_out_info_0_branchInfo_predictPC = _zz_io_out_info_0_branchInfo_predictPC;
  assign io_out_info_0_branchInfo_predictResult = _zz_io_out_info_0_branchInfo_predictResult;
  assign io_out_info_0_exceptionInfo_exception = _zz_io_out_info_0_exceptionInfo_exception;
  assign io_out_info_0_exceptionInfo_eCode = _zz_io_out_info_0_exceptionInfo_eCode;
  assign io_out_info_0_exceptionInfo_eSubCode = _zz_io_out_info_0_exceptionInfo_eSubCode;
  assign io_out_info_0_pc = _zz_io_out_info_0_pc;
  assign _zz_io_out_dispatchInfo_0_ard_1 = _zz_io_out_info_0_inst[4 : 0];
  assign _zz_when_InstrQueue_l119 = _zz_io_out_info_0_inst[9 : 5];
  assign _zz_io_out_dispatchInfo_0_asrc_1_1 = _zz_io_out_info_0_inst[14 : 10];
  assign _zz_io_out_dispatchInfo_0_ard_2 = 1'b0;
  always @(*) begin
    _zz_io_out_dispatchInfo_0_ard = {4'd0, _zz_io_out_dispatchInfo_0_ard_2};
    casez(_zz_io_out_info_0_inst)
      32'b0000000000000000011000?????00000 : begin
        _zz_io_out_dispatchInfo_0_ard = _zz_when_InstrQueue_l119;
      end
      32'b000000000000000001100000000?????, 32'b000000000000000001100100000????? : begin
        _zz_io_out_dispatchInfo_0_ard = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b00000000000100000???????????????, 32'b00000000000100010???????????????, 32'b00000000000100100???????????????, 32'b00000000000100101???????????????, 32'b00000000000101000???????????????, 32'b00000000000101001???????????????, 32'b00000000000101010???????????????, 32'b00000000000101011???????????????, 32'b00000000000101110???????????????, 32'b00000000000101111???????????????, 32'b00000000000110000??????????????? : begin
        _zz_io_out_dispatchInfo_0_ard = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b0000001010??????????????????????, 32'b0000001000??????????????????????, 32'b0000001001??????????????????????, 32'b0000001101??????????????????????, 32'b0000001110??????????????????????, 32'b0000001111??????????????????????, 32'b00000000010000001???????????????, 32'b00000000010001001???????????????, 32'b00000000010010001???????????????, 32'b010011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_0_ard = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b00000000001010100???????????????, 32'b00000000001010110???????????????, 32'b00000110010010000011100000000000, 32'b00000110010010001???????????????, 32'b010100?????????????????????????? : begin
      end
      32'b0001010?????????????????????????, 32'b0001110????????????????????????? : begin
        _zz_io_out_dispatchInfo_0_ard = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b010101?????????????????????????? : begin
        _zz_io_out_dispatchInfo_0_ard = {4'd0, _zz__zz_io_out_dispatchInfo_0_ard};
      end
      32'b010110??????????????????????????, 32'b010111??????????????????????????, 32'b011000??????????????????????????, 32'b011001??????????????????????????, 32'b011010??????????????????????????, 32'b011011?????????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
        _zz_io_out_dispatchInfo_0_ard = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b00000000000111000???????????????, 32'b00000000000111001???????????????, 32'b00000000000111010??????????????? : begin
        _zz_io_out_dispatchInfo_0_ard = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b00000000001000000???????????????, 32'b00000000001000001???????????????, 32'b00000000001000010???????????????, 32'b00000000001000011??????????????? : begin
        _zz_io_out_dispatchInfo_0_ard = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b00100000????????????????????????, 32'b0010100000??????????????????????, 32'b0010101000??????????????????????, 32'b0010100001??????????????????????, 32'b0010101001?????????????????????? : begin
        _zz_io_out_dispatchInfo_0_ard = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b0000011000??????????????????????, 32'b00000110010010011???????????????, 32'b0010101011?????????????????????? : begin
      end
      32'b00000110010010000010100000000000, 32'b00000110010010000010110000000000, 32'b00000110010010000011000000000000, 32'b00000110010010000011010000000000, 32'b00111000011100100???????????????, 32'b00111000011100101??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b00100001???????????????????????? : begin
        _zz_io_out_dispatchInfo_0_ard = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b0010100100??????????????????????, 32'b0010100101??????????????????????, 32'b0010100110?????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_out_dispatchInfo_0_asrc_0 = {4'd0, _zz_io_out_dispatchInfo_0_ard_2};
    casez(_zz_io_out_info_0_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000?????, 32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000???????????????, 32'b00000000000100010???????????????, 32'b00000000000100100???????????????, 32'b00000000000100101???????????????, 32'b00000000000101000???????????????, 32'b00000000000101001???????????????, 32'b00000000000101010???????????????, 32'b00000000000101011???????????????, 32'b00000000000101110???????????????, 32'b00000000000101111???????????????, 32'b00000000000110000??????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_0 = _zz_when_InstrQueue_l119;
      end
      32'b0000001010??????????????????????, 32'b0000001000??????????????????????, 32'b0000001001??????????????????????, 32'b0000001101??????????????????????, 32'b0000001110??????????????????????, 32'b0000001111??????????????????????, 32'b00000000010000001???????????????, 32'b00000000010001001???????????????, 32'b00000000010010001???????????????, 32'b010011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_0 = _zz_when_InstrQueue_l119;
      end
      32'b00000000001010100???????????????, 32'b00000000001010110???????????????, 32'b00000110010010000011100000000000, 32'b00000110010010001???????????????, 32'b010100?????????????????????????? : begin
      end
      32'b0001010?????????????????????????, 32'b0001110????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110??????????????????????????, 32'b010111??????????????????????????, 32'b011000??????????????????????????, 32'b011001??????????????????????????, 32'b011010??????????????????????????, 32'b011011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_0 = _zz_when_InstrQueue_l119;
      end
      32'b00000100???????????????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_0 = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b00000000000111000???????????????, 32'b00000000000111001???????????????, 32'b00000000000111010??????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_0 = _zz_when_InstrQueue_l119;
      end
      32'b00000000001000000???????????????, 32'b00000000001000001???????????????, 32'b00000000001000010???????????????, 32'b00000000001000011??????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_0 = _zz_when_InstrQueue_l119;
      end
      32'b00100000????????????????????????, 32'b0010100000??????????????????????, 32'b0010101000??????????????????????, 32'b0010100001??????????????????????, 32'b0010101001?????????????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_0 = _zz_when_InstrQueue_l119;
      end
      32'b0000011000??????????????????????, 32'b00000110010010011???????????????, 32'b0010101011?????????????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_0 = _zz_when_InstrQueue_l119;
      end
      32'b00000110010010000010100000000000, 32'b00000110010010000010110000000000, 32'b00000110010010000011000000000000, 32'b00000110010010000011010000000000, 32'b00111000011100100???????????????, 32'b00111000011100101??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_0 = _zz_when_InstrQueue_l119;
      end
      32'b00100001???????????????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_0 = _zz_when_InstrQueue_l119;
      end
      32'b0010100100??????????????????????, 32'b0010100101??????????????????????, 32'b0010100110?????????????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_0 = _zz_when_InstrQueue_l119;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_out_dispatchInfo_0_asrc_1 = {4'd0, _zz_io_out_dispatchInfo_0_ard_2};
    casez(_zz_io_out_info_0_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000?????, 32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000???????????????, 32'b00000000000100010???????????????, 32'b00000000000100100???????????????, 32'b00000000000100101???????????????, 32'b00000000000101000???????????????, 32'b00000000000101001???????????????, 32'b00000000000101010???????????????, 32'b00000000000101011???????????????, 32'b00000000000101110???????????????, 32'b00000000000101111???????????????, 32'b00000000000110000??????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_1 = _zz_io_out_dispatchInfo_0_asrc_1_1;
      end
      32'b0000001010??????????????????????, 32'b0000001000??????????????????????, 32'b0000001001??????????????????????, 32'b0000001101??????????????????????, 32'b0000001110??????????????????????, 32'b0000001111??????????????????????, 32'b00000000010000001???????????????, 32'b00000000010001001???????????????, 32'b00000000010010001???????????????, 32'b010011?????????????????????????? : begin
      end
      32'b00000000001010100???????????????, 32'b00000000001010110???????????????, 32'b00000110010010000011100000000000, 32'b00000110010010001???????????????, 32'b010100?????????????????????????? : begin
      end
      32'b0001010?????????????????????????, 32'b0001110????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110??????????????????????????, 32'b010111??????????????????????????, 32'b011000??????????????????????????, 32'b011001??????????????????????????, 32'b011010??????????????????????????, 32'b011011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_1 = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b00000100???????????????????????? : begin
        if(when_InstrQueue_l119) begin
          _zz_io_out_dispatchInfo_0_asrc_1 = _zz_when_InstrQueue_l119;
        end
      end
      32'b00000000000111000???????????????, 32'b00000000000111001???????????????, 32'b00000000000111010??????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_1 = _zz_io_out_dispatchInfo_0_asrc_1_1;
      end
      32'b00000000001000000???????????????, 32'b00000000001000001???????????????, 32'b00000000001000010???????????????, 32'b00000000001000011??????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_1 = _zz_io_out_dispatchInfo_0_asrc_1_1;
      end
      32'b00100000????????????????????????, 32'b0010100000??????????????????????, 32'b0010101000??????????????????????, 32'b0010100001??????????????????????, 32'b0010101001?????????????????????? : begin
      end
      32'b0000011000??????????????????????, 32'b00000110010010011???????????????, 32'b0010101011?????????????????????? : begin
      end
      32'b00000110010010000010100000000000, 32'b00000110010010000010110000000000, 32'b00000110010010000011000000000000, 32'b00000110010010000011010000000000, 32'b00111000011100100???????????????, 32'b00111000011100101??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_1 = _zz_io_out_dispatchInfo_0_asrc_1_1;
      end
      32'b00100001???????????????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_1 = _zz_io_out_dispatchInfo_0_ard_1;
      end
      32'b0010100100??????????????????????, 32'b0010100101??????????????????????, 32'b0010100110?????????????????????? : begin
        _zz_io_out_dispatchInfo_0_asrc_1 = _zz_io_out_dispatchInfo_0_ard_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    casez(_zz_io_out_info_0_inst)
      32'b0000000000000000011000?????00000 : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_counter;
      end
      32'b000000000000000001100000000?????, 32'b000000000000000001100100000????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_counter;
      end
      32'b00000000000100000???????????????, 32'b00000000000100010???????????????, 32'b00000000000100100???????????????, 32'b00000000000100101???????????????, 32'b00000000000101000???????????????, 32'b00000000000101001???????????????, 32'b00000000000101010???????????????, 32'b00000000000101011???????????????, 32'b00000000000101110???????????????, 32'b00000000000101111???????????????, 32'b00000000000110000??????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_alu;
      end
      32'b0000001010??????????????????????, 32'b0000001000??????????????????????, 32'b0000001001??????????????????????, 32'b0000001101??????????????????????, 32'b0000001110??????????????????????, 32'b0000001111??????????????????????, 32'b00000000010000001???????????????, 32'b00000000010001001???????????????, 32'b00000000010010001???????????????, 32'b010011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_alu;
      end
      32'b00000000001010100???????????????, 32'b00000000001010110???????????????, 32'b00000110010010000011100000000000, 32'b00000110010010001???????????????, 32'b010100?????????????????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_alu;
      end
      32'b0001010?????????????????????????, 32'b0001110????????????????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_alu;
      end
      32'b010101?????????????????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_alu;
      end
      32'b010110??????????????????????????, 32'b010111??????????????????????????, 32'b011000??????????????????????????, 32'b011001??????????????????????????, 32'b011010??????????????????????????, 32'b011011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_alu;
      end
      32'b00000100???????????????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_csr;
      end
      32'b00000000000111000???????????????, 32'b00000000000111001???????????????, 32'b00000000000111010??????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_mulu;
      end
      32'b00000000001000000???????????????, 32'b00000000001000001???????????????, 32'b00000000001000010???????????????, 32'b00000000001000011??????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_divu;
      end
      32'b00100000????????????????????????, 32'b0010100000??????????????????????, 32'b0010101000??????????????????????, 32'b0010100001??????????????????????, 32'b0010101001?????????????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_lsu;
      end
      32'b0000011000??????????????????????, 32'b00000110010010011???????????????, 32'b0010101011?????????????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_lsu;
      end
      32'b00000110010010000010100000000000, 32'b00000110010010000010110000000000, 32'b00000110010010000011000000000000, 32'b00000110010010000011010000000000, 32'b00111000011100100???????????????, 32'b00111000011100101??????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_lsu;
      end
      32'b00000110010010011??????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_lsu;
      end
      32'b00100001???????????????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_lsu;
      end
      32'b0010100100??????????????????????, 32'b0010100101??????????????????????, 32'b0010100110?????????????????????? : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_lsu;
      end
      default : begin
        _zz_io_out_dispatchInfo_0_fuType = FUType_alu;
      end
    endcase
  end

  assign when_InstrQueue_l119 = ((_zz_when_InstrQueue_l119 != 5'h00) && (_zz_when_InstrQueue_l119 != _zz_when_InstrQueue_l119_2));
  assign io_out_dispatchInfo_0_fuType = _zz_io_out_dispatchInfo_0_fuType;
  assign io_out_dispatchInfo_0_ard = _zz_io_out_dispatchInfo_0_ard;
  assign io_out_dispatchInfo_0_asrc_0 = _zz_io_out_dispatchInfo_0_asrc_0;
  assign io_out_dispatchInfo_0_asrc_1 = _zz_io_out_dispatchInfo_0_asrc_1;
  always @(*) begin
    io_out_availMask[0] = _zz_io_out_availMask;
    io_out_availMask[1] = _zz_io_out_availMask_1;
  end

  assign _zz_io_out_info_1_inst = _zz__zz_io_out_info_1_inst;
  assign io_out_info_1_inst = _zz_io_out_info_1_inst;
  assign io_out_info_1_branchInfo_predictPC = _zz_io_out_info_1_branchInfo_predictPC;
  assign io_out_info_1_branchInfo_predictResult = _zz_io_out_info_1_branchInfo_predictResult;
  assign io_out_info_1_exceptionInfo_exception = _zz_io_out_info_1_exceptionInfo_exception;
  assign io_out_info_1_exceptionInfo_eCode = _zz_io_out_info_1_exceptionInfo_eCode;
  assign io_out_info_1_exceptionInfo_eSubCode = _zz_io_out_info_1_exceptionInfo_eSubCode;
  assign io_out_info_1_pc = _zz_io_out_info_1_pc;
  assign _zz_io_out_dispatchInfo_1_ard_1 = _zz_io_out_info_1_inst[4 : 0];
  assign _zz_when_InstrQueue_l119_1 = _zz_io_out_info_1_inst[9 : 5];
  assign _zz_io_out_dispatchInfo_1_asrc_1_1 = _zz_io_out_info_1_inst[14 : 10];
  assign _zz_io_out_dispatchInfo_1_ard_2 = 1'b0;
  always @(*) begin
    _zz_io_out_dispatchInfo_1_ard = {4'd0, _zz_io_out_dispatchInfo_1_ard_2};
    casez(_zz_io_out_info_1_inst)
      32'b0000000000000000011000?????00000 : begin
        _zz_io_out_dispatchInfo_1_ard = _zz_when_InstrQueue_l119_1;
      end
      32'b000000000000000001100000000?????, 32'b000000000000000001100100000????? : begin
        _zz_io_out_dispatchInfo_1_ard = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b00000000000100000???????????????, 32'b00000000000100010???????????????, 32'b00000000000100100???????????????, 32'b00000000000100101???????????????, 32'b00000000000101000???????????????, 32'b00000000000101001???????????????, 32'b00000000000101010???????????????, 32'b00000000000101011???????????????, 32'b00000000000101110???????????????, 32'b00000000000101111???????????????, 32'b00000000000110000??????????????? : begin
        _zz_io_out_dispatchInfo_1_ard = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b0000001010??????????????????????, 32'b0000001000??????????????????????, 32'b0000001001??????????????????????, 32'b0000001101??????????????????????, 32'b0000001110??????????????????????, 32'b0000001111??????????????????????, 32'b00000000010000001???????????????, 32'b00000000010001001???????????????, 32'b00000000010010001???????????????, 32'b010011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_1_ard = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b00000000001010100???????????????, 32'b00000000001010110???????????????, 32'b00000110010010000011100000000000, 32'b00000110010010001???????????????, 32'b010100?????????????????????????? : begin
      end
      32'b0001010?????????????????????????, 32'b0001110????????????????????????? : begin
        _zz_io_out_dispatchInfo_1_ard = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b010101?????????????????????????? : begin
        _zz_io_out_dispatchInfo_1_ard = {4'd0, _zz__zz_io_out_dispatchInfo_1_ard};
      end
      32'b010110??????????????????????????, 32'b010111??????????????????????????, 32'b011000??????????????????????????, 32'b011001??????????????????????????, 32'b011010??????????????????????????, 32'b011011?????????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
        _zz_io_out_dispatchInfo_1_ard = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b00000000000111000???????????????, 32'b00000000000111001???????????????, 32'b00000000000111010??????????????? : begin
        _zz_io_out_dispatchInfo_1_ard = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b00000000001000000???????????????, 32'b00000000001000001???????????????, 32'b00000000001000010???????????????, 32'b00000000001000011??????????????? : begin
        _zz_io_out_dispatchInfo_1_ard = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b00100000????????????????????????, 32'b0010100000??????????????????????, 32'b0010101000??????????????????????, 32'b0010100001??????????????????????, 32'b0010101001?????????????????????? : begin
        _zz_io_out_dispatchInfo_1_ard = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b0000011000??????????????????????, 32'b00000110010010011???????????????, 32'b0010101011?????????????????????? : begin
      end
      32'b00000110010010000010100000000000, 32'b00000110010010000010110000000000, 32'b00000110010010000011000000000000, 32'b00000110010010000011010000000000, 32'b00111000011100100???????????????, 32'b00111000011100101??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b00100001???????????????????????? : begin
        _zz_io_out_dispatchInfo_1_ard = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b0010100100??????????????????????, 32'b0010100101??????????????????????, 32'b0010100110?????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_out_dispatchInfo_1_asrc_0 = {4'd0, _zz_io_out_dispatchInfo_1_ard_2};
    casez(_zz_io_out_info_1_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000?????, 32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000???????????????, 32'b00000000000100010???????????????, 32'b00000000000100100???????????????, 32'b00000000000100101???????????????, 32'b00000000000101000???????????????, 32'b00000000000101001???????????????, 32'b00000000000101010???????????????, 32'b00000000000101011???????????????, 32'b00000000000101110???????????????, 32'b00000000000101111???????????????, 32'b00000000000110000??????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_0 = _zz_when_InstrQueue_l119_1;
      end
      32'b0000001010??????????????????????, 32'b0000001000??????????????????????, 32'b0000001001??????????????????????, 32'b0000001101??????????????????????, 32'b0000001110??????????????????????, 32'b0000001111??????????????????????, 32'b00000000010000001???????????????, 32'b00000000010001001???????????????, 32'b00000000010010001???????????????, 32'b010011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_0 = _zz_when_InstrQueue_l119_1;
      end
      32'b00000000001010100???????????????, 32'b00000000001010110???????????????, 32'b00000110010010000011100000000000, 32'b00000110010010001???????????????, 32'b010100?????????????????????????? : begin
      end
      32'b0001010?????????????????????????, 32'b0001110????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110??????????????????????????, 32'b010111??????????????????????????, 32'b011000??????????????????????????, 32'b011001??????????????????????????, 32'b011010??????????????????????????, 32'b011011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_0 = _zz_when_InstrQueue_l119_1;
      end
      32'b00000100???????????????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_0 = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b00000000000111000???????????????, 32'b00000000000111001???????????????, 32'b00000000000111010??????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_0 = _zz_when_InstrQueue_l119_1;
      end
      32'b00000000001000000???????????????, 32'b00000000001000001???????????????, 32'b00000000001000010???????????????, 32'b00000000001000011??????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_0 = _zz_when_InstrQueue_l119_1;
      end
      32'b00100000????????????????????????, 32'b0010100000??????????????????????, 32'b0010101000??????????????????????, 32'b0010100001??????????????????????, 32'b0010101001?????????????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_0 = _zz_when_InstrQueue_l119_1;
      end
      32'b0000011000??????????????????????, 32'b00000110010010011???????????????, 32'b0010101011?????????????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_0 = _zz_when_InstrQueue_l119_1;
      end
      32'b00000110010010000010100000000000, 32'b00000110010010000010110000000000, 32'b00000110010010000011000000000000, 32'b00000110010010000011010000000000, 32'b00111000011100100???????????????, 32'b00111000011100101??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_0 = _zz_when_InstrQueue_l119_1;
      end
      32'b00100001???????????????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_0 = _zz_when_InstrQueue_l119_1;
      end
      32'b0010100100??????????????????????, 32'b0010100101??????????????????????, 32'b0010100110?????????????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_0 = _zz_when_InstrQueue_l119_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_out_dispatchInfo_1_asrc_1 = {4'd0, _zz_io_out_dispatchInfo_1_ard_2};
    casez(_zz_io_out_info_1_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000?????, 32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000???????????????, 32'b00000000000100010???????????????, 32'b00000000000100100???????????????, 32'b00000000000100101???????????????, 32'b00000000000101000???????????????, 32'b00000000000101001???????????????, 32'b00000000000101010???????????????, 32'b00000000000101011???????????????, 32'b00000000000101110???????????????, 32'b00000000000101111???????????????, 32'b00000000000110000??????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_1 = _zz_io_out_dispatchInfo_1_asrc_1_1;
      end
      32'b0000001010??????????????????????, 32'b0000001000??????????????????????, 32'b0000001001??????????????????????, 32'b0000001101??????????????????????, 32'b0000001110??????????????????????, 32'b0000001111??????????????????????, 32'b00000000010000001???????????????, 32'b00000000010001001???????????????, 32'b00000000010010001???????????????, 32'b010011?????????????????????????? : begin
      end
      32'b00000000001010100???????????????, 32'b00000000001010110???????????????, 32'b00000110010010000011100000000000, 32'b00000110010010001???????????????, 32'b010100?????????????????????????? : begin
      end
      32'b0001010?????????????????????????, 32'b0001110????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110??????????????????????????, 32'b010111??????????????????????????, 32'b011000??????????????????????????, 32'b011001??????????????????????????, 32'b011010??????????????????????????, 32'b011011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_1 = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b00000100???????????????????????? : begin
        if(when_InstrQueue_l119_1) begin
          _zz_io_out_dispatchInfo_1_asrc_1 = _zz_when_InstrQueue_l119_1;
        end
      end
      32'b00000000000111000???????????????, 32'b00000000000111001???????????????, 32'b00000000000111010??????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_1 = _zz_io_out_dispatchInfo_1_asrc_1_1;
      end
      32'b00000000001000000???????????????, 32'b00000000001000001???????????????, 32'b00000000001000010???????????????, 32'b00000000001000011??????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_1 = _zz_io_out_dispatchInfo_1_asrc_1_1;
      end
      32'b00100000????????????????????????, 32'b0010100000??????????????????????, 32'b0010101000??????????????????????, 32'b0010100001??????????????????????, 32'b0010101001?????????????????????? : begin
      end
      32'b0000011000??????????????????????, 32'b00000110010010011???????????????, 32'b0010101011?????????????????????? : begin
      end
      32'b00000110010010000010100000000000, 32'b00000110010010000010110000000000, 32'b00000110010010000011000000000000, 32'b00000110010010000011010000000000, 32'b00111000011100100???????????????, 32'b00111000011100101??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_1 = _zz_io_out_dispatchInfo_1_asrc_1_1;
      end
      32'b00100001???????????????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_1 = _zz_io_out_dispatchInfo_1_ard_1;
      end
      32'b0010100100??????????????????????, 32'b0010100101??????????????????????, 32'b0010100110?????????????????????? : begin
        _zz_io_out_dispatchInfo_1_asrc_1 = _zz_io_out_dispatchInfo_1_ard_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    casez(_zz_io_out_info_1_inst)
      32'b0000000000000000011000?????00000 : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_counter;
      end
      32'b000000000000000001100000000?????, 32'b000000000000000001100100000????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_counter;
      end
      32'b00000000000100000???????????????, 32'b00000000000100010???????????????, 32'b00000000000100100???????????????, 32'b00000000000100101???????????????, 32'b00000000000101000???????????????, 32'b00000000000101001???????????????, 32'b00000000000101010???????????????, 32'b00000000000101011???????????????, 32'b00000000000101110???????????????, 32'b00000000000101111???????????????, 32'b00000000000110000??????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_alu;
      end
      32'b0000001010??????????????????????, 32'b0000001000??????????????????????, 32'b0000001001??????????????????????, 32'b0000001101??????????????????????, 32'b0000001110??????????????????????, 32'b0000001111??????????????????????, 32'b00000000010000001???????????????, 32'b00000000010001001???????????????, 32'b00000000010010001???????????????, 32'b010011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_alu;
      end
      32'b00000000001010100???????????????, 32'b00000000001010110???????????????, 32'b00000110010010000011100000000000, 32'b00000110010010001???????????????, 32'b010100?????????????????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_alu;
      end
      32'b0001010?????????????????????????, 32'b0001110????????????????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_alu;
      end
      32'b010101?????????????????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_alu;
      end
      32'b010110??????????????????????????, 32'b010111??????????????????????????, 32'b011000??????????????????????????, 32'b011001??????????????????????????, 32'b011010??????????????????????????, 32'b011011?????????????????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_alu;
      end
      32'b00000100???????????????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_csr;
      end
      32'b00000000000111000???????????????, 32'b00000000000111001???????????????, 32'b00000000000111010??????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_mulu;
      end
      32'b00000000001000000???????????????, 32'b00000000001000001???????????????, 32'b00000000001000010???????????????, 32'b00000000001000011??????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_divu;
      end
      32'b00100000????????????????????????, 32'b0010100000??????????????????????, 32'b0010101000??????????????????????, 32'b0010100001??????????????????????, 32'b0010101001?????????????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_lsu;
      end
      32'b0000011000??????????????????????, 32'b00000110010010011???????????????, 32'b0010101011?????????????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_lsu;
      end
      32'b00000110010010000010100000000000, 32'b00000110010010000010110000000000, 32'b00000110010010000011000000000000, 32'b00000110010010000011010000000000, 32'b00111000011100100???????????????, 32'b00111000011100101??????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_lsu;
      end
      32'b00000110010010011??????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_lsu;
      end
      32'b00100001???????????????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_lsu;
      end
      32'b0010100100??????????????????????, 32'b0010100101??????????????????????, 32'b0010100110?????????????????????? : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_lsu;
      end
      default : begin
        _zz_io_out_dispatchInfo_1_fuType = FUType_alu;
      end
    endcase
  end

  assign when_InstrQueue_l119_1 = ((_zz_when_InstrQueue_l119_1 != 5'h00) && (_zz_when_InstrQueue_l119_1 != _zz_when_InstrQueue_l119_1_1));
  assign io_out_dispatchInfo_1_fuType = _zz_io_out_dispatchInfo_1_fuType;
  assign io_out_dispatchInfo_1_ard = _zz_io_out_dispatchInfo_1_ard;
  assign io_out_dispatchInfo_1_asrc_0 = _zz_io_out_dispatchInfo_1_asrc_0;
  assign io_out_dispatchInfo_1_asrc_1 = _zz_io_out_dispatchInfo_1_asrc_1;
  always @(*) begin
    _zz_valid_0[0] = ((tail_0 == 3'b000) && io_in_allowMask[0]);
    _zz_valid_0[1] = ((tail_1 == 3'b000) && io_in_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_0_1[0] = ((head_0 == 3'b000) && io_out_allowMask[0]);
    _zz_valid_0_1[1] = ((head_1 == 3'b000) && io_out_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_1[0] = ((tail_0 == 3'b001) && io_in_allowMask[0]);
    _zz_valid_1[1] = ((tail_1 == 3'b001) && io_in_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_1_1[0] = ((head_0 == 3'b001) && io_out_allowMask[0]);
    _zz_valid_1_1[1] = ((head_1 == 3'b001) && io_out_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_2[0] = ((tail_0 == 3'b010) && io_in_allowMask[0]);
    _zz_valid_2[1] = ((tail_1 == 3'b010) && io_in_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_2_1[0] = ((head_0 == 3'b010) && io_out_allowMask[0]);
    _zz_valid_2_1[1] = ((head_1 == 3'b010) && io_out_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_3[0] = ((tail_0 == 3'b011) && io_in_allowMask[0]);
    _zz_valid_3[1] = ((tail_1 == 3'b011) && io_in_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_3_1[0] = ((head_0 == 3'b011) && io_out_allowMask[0]);
    _zz_valid_3_1[1] = ((head_1 == 3'b011) && io_out_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_4[0] = ((tail_0 == 3'b100) && io_in_allowMask[0]);
    _zz_valid_4[1] = ((tail_1 == 3'b100) && io_in_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_4_1[0] = ((head_0 == 3'b100) && io_out_allowMask[0]);
    _zz_valid_4_1[1] = ((head_1 == 3'b100) && io_out_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_5[0] = ((tail_0 == 3'b101) && io_in_allowMask[0]);
    _zz_valid_5[1] = ((tail_1 == 3'b101) && io_in_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_5_1[0] = ((head_0 == 3'b101) && io_out_allowMask[0]);
    _zz_valid_5_1[1] = ((head_1 == 3'b101) && io_out_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_6[0] = ((tail_0 == 3'b110) && io_in_allowMask[0]);
    _zz_valid_6[1] = ((tail_1 == 3'b110) && io_in_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_6_1[0] = ((head_0 == 3'b110) && io_out_allowMask[0]);
    _zz_valid_6_1[1] = ((head_1 == 3'b110) && io_out_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_7[0] = ((tail_0 == 3'b111) && io_in_allowMask[0]);
    _zz_valid_7[1] = ((tail_1 == 3'b111) && io_in_allowMask[1]);
  end

  always @(*) begin
    _zz_valid_7_1[0] = ((head_0 == 3'b111) && io_out_allowMask[0]);
    _zz_valid_7_1[1] = ((head_1 == 3'b111) && io_out_allowMask[1]);
  end

  always @(posedge aclk) begin
    if(!cpuClockingArea_areaFlushReset_newReset) begin
      valid_0 <= 1'b0;
      valid_1 <= 1'b0;
      valid_2 <= 1'b0;
      valid_3 <= 1'b0;
      valid_4 <= 1'b0;
      valid_5 <= 1'b0;
      valid_6 <= 1'b0;
      valid_7 <= 1'b0;
      head_0 <= 3'b000;
      head_1 <= 3'b001;
      tail_0 <= 3'b000;
      tail_1 <= 3'b001;
    end else begin
      tail_0 <= (tail_0 + _zz_tail_0);
      tail_1 <= (tail_1 + _zz_tail_1);
      head_0 <= (head_0 + _zz_head_0);
      head_1 <= (head_1 + _zz_head_1);
      valid_0 <= ((|_zz_valid_0_1) ? 1'b0 : (valid_0 || (|_zz_valid_0)));
      valid_1 <= ((|_zz_valid_1_1) ? 1'b0 : (valid_1 || (|_zz_valid_1)));
      valid_2 <= ((|_zz_valid_2_1) ? 1'b0 : (valid_2 || (|_zz_valid_2)));
      valid_3 <= ((|_zz_valid_3_1) ? 1'b0 : (valid_3 || (|_zz_valid_3)));
      valid_4 <= ((|_zz_valid_4_1) ? 1'b0 : (valid_4 || (|_zz_valid_4)));
      valid_5 <= ((|_zz_valid_5_1) ? 1'b0 : (valid_5 || (|_zz_valid_5)));
      valid_6 <= ((|_zz_valid_6_1) ? 1'b0 : (valid_6 || (|_zz_valid_6)));
      valid_7 <= ((|_zz_valid_7_1) ? 1'b0 : (valid_7 || (|_zz_valid_7)));
    end
  end

  always @(posedge aclk) begin
    if(when_InstrQueue_l33) begin
      if(_zz_2) begin
        queue_0_inst <= io_in_info_0_inst;
      end
      if(_zz_3) begin
        queue_1_inst <= io_in_info_0_inst;
      end
      if(_zz_4) begin
        queue_2_inst <= io_in_info_0_inst;
      end
      if(_zz_5) begin
        queue_3_inst <= io_in_info_0_inst;
      end
      if(_zz_6) begin
        queue_4_inst <= io_in_info_0_inst;
      end
      if(_zz_7) begin
        queue_5_inst <= io_in_info_0_inst;
      end
      if(_zz_8) begin
        queue_6_inst <= io_in_info_0_inst;
      end
      if(_zz_9) begin
        queue_7_inst <= io_in_info_0_inst;
      end
      if(_zz_2) begin
        queue_0_branchInfo_predictPC <= io_in_info_0_branchInfo_predictPC;
      end
      if(_zz_3) begin
        queue_1_branchInfo_predictPC <= io_in_info_0_branchInfo_predictPC;
      end
      if(_zz_4) begin
        queue_2_branchInfo_predictPC <= io_in_info_0_branchInfo_predictPC;
      end
      if(_zz_5) begin
        queue_3_branchInfo_predictPC <= io_in_info_0_branchInfo_predictPC;
      end
      if(_zz_6) begin
        queue_4_branchInfo_predictPC <= io_in_info_0_branchInfo_predictPC;
      end
      if(_zz_7) begin
        queue_5_branchInfo_predictPC <= io_in_info_0_branchInfo_predictPC;
      end
      if(_zz_8) begin
        queue_6_branchInfo_predictPC <= io_in_info_0_branchInfo_predictPC;
      end
      if(_zz_9) begin
        queue_7_branchInfo_predictPC <= io_in_info_0_branchInfo_predictPC;
      end
      if(_zz_2) begin
        queue_0_branchInfo_predictResult <= io_in_info_0_branchInfo_predictResult;
      end
      if(_zz_3) begin
        queue_1_branchInfo_predictResult <= io_in_info_0_branchInfo_predictResult;
      end
      if(_zz_4) begin
        queue_2_branchInfo_predictResult <= io_in_info_0_branchInfo_predictResult;
      end
      if(_zz_5) begin
        queue_3_branchInfo_predictResult <= io_in_info_0_branchInfo_predictResult;
      end
      if(_zz_6) begin
        queue_4_branchInfo_predictResult <= io_in_info_0_branchInfo_predictResult;
      end
      if(_zz_7) begin
        queue_5_branchInfo_predictResult <= io_in_info_0_branchInfo_predictResult;
      end
      if(_zz_8) begin
        queue_6_branchInfo_predictResult <= io_in_info_0_branchInfo_predictResult;
      end
      if(_zz_9) begin
        queue_7_branchInfo_predictResult <= io_in_info_0_branchInfo_predictResult;
      end
      if(_zz_2) begin
        queue_0_exceptionInfo_exception <= io_in_info_0_exceptionInfo_exception;
      end
      if(_zz_3) begin
        queue_1_exceptionInfo_exception <= io_in_info_0_exceptionInfo_exception;
      end
      if(_zz_4) begin
        queue_2_exceptionInfo_exception <= io_in_info_0_exceptionInfo_exception;
      end
      if(_zz_5) begin
        queue_3_exceptionInfo_exception <= io_in_info_0_exceptionInfo_exception;
      end
      if(_zz_6) begin
        queue_4_exceptionInfo_exception <= io_in_info_0_exceptionInfo_exception;
      end
      if(_zz_7) begin
        queue_5_exceptionInfo_exception <= io_in_info_0_exceptionInfo_exception;
      end
      if(_zz_8) begin
        queue_6_exceptionInfo_exception <= io_in_info_0_exceptionInfo_exception;
      end
      if(_zz_9) begin
        queue_7_exceptionInfo_exception <= io_in_info_0_exceptionInfo_exception;
      end
      if(_zz_2) begin
        queue_0_exceptionInfo_eCode <= io_in_info_0_exceptionInfo_eCode;
      end
      if(_zz_3) begin
        queue_1_exceptionInfo_eCode <= io_in_info_0_exceptionInfo_eCode;
      end
      if(_zz_4) begin
        queue_2_exceptionInfo_eCode <= io_in_info_0_exceptionInfo_eCode;
      end
      if(_zz_5) begin
        queue_3_exceptionInfo_eCode <= io_in_info_0_exceptionInfo_eCode;
      end
      if(_zz_6) begin
        queue_4_exceptionInfo_eCode <= io_in_info_0_exceptionInfo_eCode;
      end
      if(_zz_7) begin
        queue_5_exceptionInfo_eCode <= io_in_info_0_exceptionInfo_eCode;
      end
      if(_zz_8) begin
        queue_6_exceptionInfo_eCode <= io_in_info_0_exceptionInfo_eCode;
      end
      if(_zz_9) begin
        queue_7_exceptionInfo_eCode <= io_in_info_0_exceptionInfo_eCode;
      end
      if(_zz_2) begin
        queue_0_exceptionInfo_eSubCode <= io_in_info_0_exceptionInfo_eSubCode;
      end
      if(_zz_3) begin
        queue_1_exceptionInfo_eSubCode <= io_in_info_0_exceptionInfo_eSubCode;
      end
      if(_zz_4) begin
        queue_2_exceptionInfo_eSubCode <= io_in_info_0_exceptionInfo_eSubCode;
      end
      if(_zz_5) begin
        queue_3_exceptionInfo_eSubCode <= io_in_info_0_exceptionInfo_eSubCode;
      end
      if(_zz_6) begin
        queue_4_exceptionInfo_eSubCode <= io_in_info_0_exceptionInfo_eSubCode;
      end
      if(_zz_7) begin
        queue_5_exceptionInfo_eSubCode <= io_in_info_0_exceptionInfo_eSubCode;
      end
      if(_zz_8) begin
        queue_6_exceptionInfo_eSubCode <= io_in_info_0_exceptionInfo_eSubCode;
      end
      if(_zz_9) begin
        queue_7_exceptionInfo_eSubCode <= io_in_info_0_exceptionInfo_eSubCode;
      end
      if(_zz_2) begin
        queue_0_pc <= io_in_info_0_pc;
      end
      if(_zz_3) begin
        queue_1_pc <= io_in_info_0_pc;
      end
      if(_zz_4) begin
        queue_2_pc <= io_in_info_0_pc;
      end
      if(_zz_5) begin
        queue_3_pc <= io_in_info_0_pc;
      end
      if(_zz_6) begin
        queue_4_pc <= io_in_info_0_pc;
      end
      if(_zz_7) begin
        queue_5_pc <= io_in_info_0_pc;
      end
      if(_zz_8) begin
        queue_6_pc <= io_in_info_0_pc;
      end
      if(_zz_9) begin
        queue_7_pc <= io_in_info_0_pc;
      end
    end
    if(when_InstrQueue_l33_1) begin
      if(_zz_11) begin
        queue_0_inst <= io_in_info_1_inst;
      end
      if(_zz_12) begin
        queue_1_inst <= io_in_info_1_inst;
      end
      if(_zz_13) begin
        queue_2_inst <= io_in_info_1_inst;
      end
      if(_zz_14) begin
        queue_3_inst <= io_in_info_1_inst;
      end
      if(_zz_15) begin
        queue_4_inst <= io_in_info_1_inst;
      end
      if(_zz_16) begin
        queue_5_inst <= io_in_info_1_inst;
      end
      if(_zz_17) begin
        queue_6_inst <= io_in_info_1_inst;
      end
      if(_zz_18) begin
        queue_7_inst <= io_in_info_1_inst;
      end
      if(_zz_11) begin
        queue_0_branchInfo_predictPC <= io_in_info_1_branchInfo_predictPC;
      end
      if(_zz_12) begin
        queue_1_branchInfo_predictPC <= io_in_info_1_branchInfo_predictPC;
      end
      if(_zz_13) begin
        queue_2_branchInfo_predictPC <= io_in_info_1_branchInfo_predictPC;
      end
      if(_zz_14) begin
        queue_3_branchInfo_predictPC <= io_in_info_1_branchInfo_predictPC;
      end
      if(_zz_15) begin
        queue_4_branchInfo_predictPC <= io_in_info_1_branchInfo_predictPC;
      end
      if(_zz_16) begin
        queue_5_branchInfo_predictPC <= io_in_info_1_branchInfo_predictPC;
      end
      if(_zz_17) begin
        queue_6_branchInfo_predictPC <= io_in_info_1_branchInfo_predictPC;
      end
      if(_zz_18) begin
        queue_7_branchInfo_predictPC <= io_in_info_1_branchInfo_predictPC;
      end
      if(_zz_11) begin
        queue_0_branchInfo_predictResult <= io_in_info_1_branchInfo_predictResult;
      end
      if(_zz_12) begin
        queue_1_branchInfo_predictResult <= io_in_info_1_branchInfo_predictResult;
      end
      if(_zz_13) begin
        queue_2_branchInfo_predictResult <= io_in_info_1_branchInfo_predictResult;
      end
      if(_zz_14) begin
        queue_3_branchInfo_predictResult <= io_in_info_1_branchInfo_predictResult;
      end
      if(_zz_15) begin
        queue_4_branchInfo_predictResult <= io_in_info_1_branchInfo_predictResult;
      end
      if(_zz_16) begin
        queue_5_branchInfo_predictResult <= io_in_info_1_branchInfo_predictResult;
      end
      if(_zz_17) begin
        queue_6_branchInfo_predictResult <= io_in_info_1_branchInfo_predictResult;
      end
      if(_zz_18) begin
        queue_7_branchInfo_predictResult <= io_in_info_1_branchInfo_predictResult;
      end
      if(_zz_11) begin
        queue_0_exceptionInfo_exception <= io_in_info_1_exceptionInfo_exception;
      end
      if(_zz_12) begin
        queue_1_exceptionInfo_exception <= io_in_info_1_exceptionInfo_exception;
      end
      if(_zz_13) begin
        queue_2_exceptionInfo_exception <= io_in_info_1_exceptionInfo_exception;
      end
      if(_zz_14) begin
        queue_3_exceptionInfo_exception <= io_in_info_1_exceptionInfo_exception;
      end
      if(_zz_15) begin
        queue_4_exceptionInfo_exception <= io_in_info_1_exceptionInfo_exception;
      end
      if(_zz_16) begin
        queue_5_exceptionInfo_exception <= io_in_info_1_exceptionInfo_exception;
      end
      if(_zz_17) begin
        queue_6_exceptionInfo_exception <= io_in_info_1_exceptionInfo_exception;
      end
      if(_zz_18) begin
        queue_7_exceptionInfo_exception <= io_in_info_1_exceptionInfo_exception;
      end
      if(_zz_11) begin
        queue_0_exceptionInfo_eCode <= io_in_info_1_exceptionInfo_eCode;
      end
      if(_zz_12) begin
        queue_1_exceptionInfo_eCode <= io_in_info_1_exceptionInfo_eCode;
      end
      if(_zz_13) begin
        queue_2_exceptionInfo_eCode <= io_in_info_1_exceptionInfo_eCode;
      end
      if(_zz_14) begin
        queue_3_exceptionInfo_eCode <= io_in_info_1_exceptionInfo_eCode;
      end
      if(_zz_15) begin
        queue_4_exceptionInfo_eCode <= io_in_info_1_exceptionInfo_eCode;
      end
      if(_zz_16) begin
        queue_5_exceptionInfo_eCode <= io_in_info_1_exceptionInfo_eCode;
      end
      if(_zz_17) begin
        queue_6_exceptionInfo_eCode <= io_in_info_1_exceptionInfo_eCode;
      end
      if(_zz_18) begin
        queue_7_exceptionInfo_eCode <= io_in_info_1_exceptionInfo_eCode;
      end
      if(_zz_11) begin
        queue_0_exceptionInfo_eSubCode <= io_in_info_1_exceptionInfo_eSubCode;
      end
      if(_zz_12) begin
        queue_1_exceptionInfo_eSubCode <= io_in_info_1_exceptionInfo_eSubCode;
      end
      if(_zz_13) begin
        queue_2_exceptionInfo_eSubCode <= io_in_info_1_exceptionInfo_eSubCode;
      end
      if(_zz_14) begin
        queue_3_exceptionInfo_eSubCode <= io_in_info_1_exceptionInfo_eSubCode;
      end
      if(_zz_15) begin
        queue_4_exceptionInfo_eSubCode <= io_in_info_1_exceptionInfo_eSubCode;
      end
      if(_zz_16) begin
        queue_5_exceptionInfo_eSubCode <= io_in_info_1_exceptionInfo_eSubCode;
      end
      if(_zz_17) begin
        queue_6_exceptionInfo_eSubCode <= io_in_info_1_exceptionInfo_eSubCode;
      end
      if(_zz_18) begin
        queue_7_exceptionInfo_eSubCode <= io_in_info_1_exceptionInfo_eSubCode;
      end
      if(_zz_11) begin
        queue_0_pc <= io_in_info_1_pc;
      end
      if(_zz_12) begin
        queue_1_pc <= io_in_info_1_pc;
      end
      if(_zz_13) begin
        queue_2_pc <= io_in_info_1_pc;
      end
      if(_zz_14) begin
        queue_3_pc <= io_in_info_1_pc;
      end
      if(_zz_15) begin
        queue_4_pc <= io_in_info_1_pc;
      end
      if(_zz_16) begin
        queue_5_pc <= io_in_info_1_pc;
      end
      if(_zz_17) begin
        queue_6_pc <= io_in_info_1_pc;
      end
      if(_zz_18) begin
        queue_7_pc <= io_in_info_1_pc;
      end
    end
  end


endmodule

module CSR (
  input  wire [7:0]    io_extInt,
  output wire          io_interrupt,
  output wire [1:0]    _zz_when_Cache_l83,
  output wire [31:0]   io_counter_id,
  output wire [63:0]   io_counter_value,
  output reg  [31:0]   io_swRead_value,
  input  wire [13:0]   io_swRead_address,
  input  wire [31:0]   io_swWrite_value,
  input  wire [13:0]   io_swWrite_address,
  input  wire          io_swWrite_wen,
  output wire [31:0]   io_llBitComm_actualAddr,
  input  wire [31:0]   io_llBitComm_toUpdateAddr,
  input  wire          io_llBitComm_wen,
  output wire          _zz_scMatchHit,
  input  wire [31:0]   io_badvICache_vaddr,
  input  wire          io_badvICache_wen,
  input  wire [4:0]    io_badvDCache_robIdx,
  input  wire [31:0]   io_badvDCache_vaddr,
  input  wire          io_badvDCache_wen,
  output wire [9:0]    io_tlbCSRInfo_asid,
  output wire [1:0]    _zz_io_iCacheReq_pageInfo_plv,
  output wire          _zz_when_TLB_l177,
  output wire          _zz_when_TLB_l177_1,
  output wire [1:0]    _zz_io_iCacheReq_pageInfo_mat,
  output wire [1:0]    _zz_io_dCacheReq_pageInfo_mat,
  output wire          _zz_when_TLB_l178,
  output wire          _zz_when_TLB_l178_1,
  output wire [1:0]    _zz_io_iCacheReq_pageInfo_mat_1,
  output wire [2:0]    _zz_io_iCacheReq_pageInfo_ppn,
  output wire [2:0]    _zz_when_TLB_l178_2,
  output wire          _zz_when_TLB_l185,
  output wire          _zz_when_TLB_l185_1,
  output wire [1:0]    _zz_io_iCacheReq_pageInfo_mat_2,
  output wire [2:0]    _zz_io_iCacheReq_pageInfo_ppn_1,
  output wire [2:0]    _zz_when_TLB_l185_2,
  output wire [5:0]    _zz_entryToFill_e,
  output wire [1:0]    _zz_io_csrWrite_asid,
  output wire [21:0]   _zz_io_swRead_value,
  output wire [5:0]    _zz_entryToFill_ps,
  output wire          _zz_io_swRead_value_1,
  output wire          _zz_entryToFill_e_1,
  output wire [18:0]   _zz_entryToFill_vppn,
  output wire          _zz_entryToFill_pp0_v,
  output wire          _zz_entryToFill_pp0_d,
  output wire [1:0]    _zz_entryToFill_pp0_plv,
  output wire [1:0]    _zz_entryToFill_pp0_mat,
  output wire          _zz_entryToFill_g,
  output wire [19:0]   _zz_entryToFill_pp0_ppn,
  output wire          _zz_entryToFill_pp1_v,
  output wire          _zz_entryToFill_pp1_d,
  output wire [1:0]    _zz_entryToFill_pp1_plv,
  output wire [1:0]    _zz_entryToFill_pp1_mat,
  output wire          _zz_entryToFill_g_1,
  output wire [19:0]   _zz_entryToFill_pp1_ppn,
  input  wire [1:0]    _zz_io_swRead_value_2,
  input  wire [21:0]   _zz_io_swRead_value_3,
  input  wire [5:0]    _zz_io_swRead_value_4,
  input  wire          _zz_io_swRead_value_5,
  input  wire          _zz_io_swRead_value_6,
  input  wire [12:0]   _zz_io_swRead_value_7,
  input  wire [18:0]   _zz_io_swRead_value_8,
  input  wire          _zz_io_swRead_value_9,
  input  wire          _zz_io_swRead_value_10,
  input  wire [1:0]    _zz_io_swRead_value_11,
  input  wire [1:0]    _zz_io_swRead_value_12,
  input  wire          _zz_io_swRead_value_13,
  input  wire          _zz_io_swRead_value_14,
  input  wire [19:0]   _zz_io_swRead_value_15,
  input  wire [3:0]    _zz_io_swRead_value_16,
  input  wire          _zz_io_swRead_value_17,
  input  wire          _zz_io_swRead_value_18,
  input  wire [1:0]    _zz_io_swRead_value_19,
  input  wire [1:0]    _zz_io_swRead_value_20,
  input  wire          _zz_io_swRead_value_21,
  input  wire          _zz_io_swRead_value_22,
  input  wire [19:0]   _zz_io_swRead_value_23,
  input  wire [3:0]    _zz_io_swRead_value_24,
  input  wire [9:0]    io_tlbCSRWrite_asid,
  input  wire          io_tlbCSRWrite_idxWen,
  input  wire          io_tlbCSRWrite_entryWen,
  input  wire          io_ctrl_llBitUpdate,
  input  wire          io_ctrl_writeCSR,
  input  wire          io_ctrl_ertn,
  input  wire          io_ctrl_normalException,
  input  wire          io_ctrl_tlbrException,
  input  wire [31:0]   io_ctrl_epc,
  input  wire [4:0]    io_ctrl_eROBIdx,
  input  wire [5:0]    io_ctrl_eCode,
  input  wire [0:0]    io_ctrl_eSubCode,
  output wire [31:0]   io_ctrl_era,
  output wire [31:0]   io_ctrl_eentry,
  output wire [31:0]   io_ctrl_tlbrentry,
  input  wire          io_flush,
  output wire [31:0]   io_diffCSRBundle_crmd,
  output wire [31:0]   io_diffCSRBundle_prmd,
  output wire [31:0]   io_diffCSRBundle_ecfg,
  output wire [31:0]   io_diffCSRBundle_estat,
  output wire [31:0]   io_diffCSRBundle_era,
  output wire [31:0]   io_diffCSRBundle_badv,
  output wire [31:0]   io_diffCSRBundle_eentry,
  output wire [31:0]   io_diffCSRBundle_tlbidx,
  output wire [31:0]   io_diffCSRBundle_tlbehi,
  output wire [31:0]   io_diffCSRBundle_tlbelo0,
  output wire [31:0]   io_diffCSRBundle_tlbelo1,
  output wire [31:0]   io_diffCSRBundle_asid,
  output wire [31:0]   io_diffCSRBundle_pgdl,
  output wire [31:0]   io_diffCSRBundle_pgdh,
  output wire [31:0]   io_diffCSRBundle_save0,
  output wire [31:0]   io_diffCSRBundle_save1,
  output wire [31:0]   io_diffCSRBundle_save2,
  output wire [31:0]   io_diffCSRBundle_save3,
  output wire [31:0]   io_diffCSRBundle_tid,
  output wire [31:0]   io_diffCSRBundle_tcfg,
  output wire [31:0]   io_diffCSRBundle_tval,
  output wire [31:0]   io_diffCSRBundle_ticlr,
  output wire [31:0]   io_diffCSRBundle_llbctl,
  output wire [31:0]   io_diffCSRBundle_tlbrentry,
  output wire [31:0]   io_diffCSRBundle_dmw0,
  output wire [31:0]   io_diffCSRBundle_dmw1,
  input  wire          aclk,
  input  wire          aresetn
);

  wire       [3:0]    _zz__zz_io_swRead_value_76;
  wire       [0:0]    _zz_io_diffCSRBundle_ticlr;
  wire       [63:0]   _zz_stableCounter_valueNext;
  wire       [0:0]    _zz_stableCounter_valueNext_1;
  wire       [31:0]   _zz__zz_io_swRead_value_112;
  wire       [31:0]   _zz__zz_io_swRead_value_112_1;
  wire       [0:0]    _zz__zz_io_swRead_value_112_2;
  wire       [31:0]   _zz_intVec;
  wire       [31:0]   _zz_intVec_1;
  wire       [31:0]   _zz__zz_io_interrupt_1;
  wire       [31:0]   _zz__zz_io_swRead_value_113;
  wire       [31:0]   _zz__zz_io_swRead_value_114;
  wire       [31:0]   _zz__zz_io_swRead_value_114_1;
  wire       [31:0]   _zz__zz_io_swRead_value_115;
  wire       [31:0]   _zz__zz_io_swRead_value_116;
  wire       [31:0]   _zz__zz_io_swRead_value_117;
  wire       [31:0]   _zz__zz_io_swRead_value_117_1;
  wire       [31:0]   _zz__zz_io_swRead_value_118;
  wire       [31:0]   _zz__zz_io_swRead_value_119;
  wire       [31:0]   _zz__zz_io_swRead_value_119_1;
  wire       [31:0]   _zz__zz_io_swRead_value_120;
  wire       [31:0]   _zz__zz_io_swRead_value_120_1;
  wire       [31:0]   _zz__zz_io_swRead_value_121;
  wire       [31:0]   _zz__zz_io_swRead_value_122;
  wire       [31:0]   _zz__zz_io_swRead_value_123;
  wire       [31:0]   _zz__zz_io_swRead_value_124;
  wire       [31:0]   _zz__zz_io_swRead_value_124_1;
  wire       [31:0]   _zz__zz_io_swRead_value_125;
  wire       [31:0]   _zz__zz_io_swRead_value_126;
  wire       [31:0]   _zz__zz_io_swRead_value_126_1;
  wire       [31:0]   _zz__zz_io_swRead_value_126_2;
  wire       [31:0]   _zz__zz_io_swRead_value_127;
  wire       [31:0]   _zz__zz_io_swRead_value_127_1;
  wire       [31:0]   _zz__zz_io_swRead_value_127_2;
  wire                _zz_when_CSR_l303;
  wire                _zz_when_CSR_l303_1;
  wire                _zz_when_CSR_l303_2;
  wire       [5:0]    _zz_when_CSR_l303_3;
  wire       [0:0]    _zz_when_CSR_l303_4;
  wire                _zz_when_CSR_l303_5;
  wire       [5:0]    _zz_when_CSR_l303_6;
  wire       [1:0]    _zz_when_CSR_l303_7;
  wire       [0:0]    _zz_when_CSR_l303_8;
  wire       [5:0]    _zz_when_CSR_l303_9;
  wire       [1:0]    _zz_when_CSR_l303_10;
  wire       [5:0]    _zz_when_CSR_l303_11;
  wire       [2:0]    _zz_when_CSR_l303_12;
  wire       [5:0]    _zz_when_CSR_l303_13;
  wire       [2:0]    _zz_when_CSR_l303_14;
  wire       [5:0]    _zz_when_CSR_l313;
  wire       [3:0]    _zz_when_CSR_l313_1;
  wire       [5:0]    _zz_when_CSR_l313_2;
  wire       [3:0]    _zz_when_CSR_l313_3;
  reg        [1:0]    _zz_io_swRead_value_25;
  reg                 _zz_io_interrupt;
  reg                 _zz_io_swRead_value_26;
  reg                 _zz_io_swRead_value_27;
  reg        [1:0]    _zz_io_swRead_value_28;
  reg        [1:0]    _zz_io_swRead_value_29;
  reg        [22:0]   _zz_io_swRead_value_30;
  reg        [1:0]    _zz_io_swRead_value_31;
  reg                 _zz_io_swRead_value_32;
  reg        [28:0]   _zz_io_swRead_value_33;
  reg        [9:0]    _zz_io_swRead_value_34;
  reg                 _zz_io_swRead_value_35;
  reg        [1:0]    _zz_io_swRead_value_36;
  reg        [18:0]   _zz_io_swRead_value_37;
  reg        [1:0]    _zz_io_swRead_value_38;
  reg        [7:0]    _zz_io_swRead_value_39;
  reg                 _zz_io_swRead_value_40;
  reg                 _zz_io_swRead_value_41;
  reg                 _zz_io_swRead_value_42;
  reg        [2:0]    _zz_io_swRead_value_43;
  reg        [5:0]    _zz_io_swRead_value_44;
  reg        [8:0]    _zz_io_swRead_value_45;
  reg                 _zz_io_swRead_value_46;
  reg        [31:0]   _zz_io_swRead_value_47;
  reg        [31:0]   _zz_io_swRead_value_48;
  reg        [5:0]    _zz_io_swRead_value_49;
  reg        [25:0]   _zz_io_swRead_value_50;
  reg        [1:0]    _zz_io_swRead_value_51;
  reg        [21:0]   _zz_io_swRead_value_52;
  reg        [5:0]    _zz_io_swRead_value_53;
  reg                 _zz_io_swRead_value_54;
  reg                 _zz_io_swRead_value_55;
  reg        [12:0]   _zz_io_swRead_value_56;
  reg        [18:0]   _zz_io_swRead_value_57;
  reg                 _zz_io_swRead_value_58;
  reg                 _zz_io_swRead_value_59;
  reg        [1:0]    _zz_io_swRead_value_60;
  reg        [1:0]    _zz_io_swRead_value_61;
  reg                 _zz_io_swRead_value_62;
  reg                 _zz_io_swRead_value_63;
  reg        [19:0]   _zz_io_swRead_value_64;
  reg        [3:0]    _zz_io_swRead_value_65;
  reg                 _zz_io_swRead_value_66;
  reg                 _zz_io_swRead_value_67;
  reg        [1:0]    _zz_io_swRead_value_68;
  reg        [1:0]    _zz_io_swRead_value_69;
  reg                 _zz_io_swRead_value_70;
  reg                 _zz_io_swRead_value_71;
  reg        [19:0]   _zz_io_swRead_value_72;
  reg        [3:0]    _zz_io_swRead_value_73;
  reg        [9:0]    _zz_io_swRead_value_74;
  reg        [5:0]    _zz_io_swRead_value_75;
  reg        [7:0]    _zz_io_swRead_value_76;
  reg        [7:0]    _zz_io_swRead_value_77;
  reg        [11:0]   _zz_io_swRead_value_78;
  reg        [19:0]   _zz_io_swRead_value_79;
  reg        [11:0]   _zz_io_swRead_value_80;
  reg        [19:0]   _zz_io_swRead_value_81;
  reg        [31:0]   _zz_io_swRead_value_82;
  reg        [31:0]   _zz_io_swRead_value_83;
  reg        [31:0]   _zz_io_swRead_value_84;
  reg        [31:0]   _zz_io_swRead_value_85;
  reg        [31:0]   _zz_io_counter_id;
  reg                 _zz_io_swRead_value_86;
  reg                 _zz_io_swRead_value_87;
  reg        [29:0]   _zz_io_swRead_value_88;
  reg        [31:0]   _zz_io_swRead_value_89;
  reg                 ticlr;
  reg                 _zz_io_swRead_value_90;
  reg                 _zz_io_swRead_value_91;
  reg                 _zz_io_swRead_value_92;
  reg        [28:0]   _zz_io_swRead_value_93;
  reg        [5:0]    _zz_io_swRead_value_94;
  reg        [25:0]   _zz_io_swRead_value_95;
  reg                 _zz_io_swRead_value_96;
  reg        [1:0]    _zz_io_swRead_value_97;
  reg                 _zz_io_swRead_value_98;
  reg        [1:0]    _zz_io_swRead_value_99;
  reg        [18:0]   _zz_io_swRead_value_100;
  reg        [2:0]    _zz_io_swRead_value_101;
  reg                 _zz_io_swRead_value_102;
  reg        [2:0]    _zz_io_swRead_value_103;
  reg                 _zz_io_swRead_value_104;
  reg        [1:0]    _zz_io_swRead_value_105;
  reg                 _zz_io_swRead_value_106;
  reg        [1:0]    _zz_io_swRead_value_107;
  reg        [18:0]   _zz_io_swRead_value_108;
  reg        [2:0]    _zz_io_swRead_value_109;
  reg                 _zz_io_swRead_value_110;
  reg        [2:0]    _zz_io_swRead_value_111;
  reg                 stableCounter_willIncrement;
  wire                stableCounter_willClear;
  reg        [63:0]   stableCounter_valueNext;
  reg        [63:0]   stableCounter_value;
  wire                stableCounter_willOverflowIfInc;
  wire                stableCounter_willOverflow;
  reg        [31:0]   _zz_io_swRead_value_112;
  wire                timeUp;
  wire                when_CSR_l116;
  wire                when_CSR_l117;
  wire       [15:0]   intVec;
  reg        [31:0]   csrWriteBuffer_value;
  reg        [13:0]   csrWriteBuffer_address;
  reg                 csrWriteBufferLock;
  wire                when_CSR_l139;
  wire                when_CSR_l143;
  reg        [31:0]   llAddr;
  reg        [31:0]   llbUpdateBuffer;
  reg                 llbUpdateBufferLock;
  wire                when_CSR_l156;
  wire                when_CSR_l159;
  reg        [31:0]   badvICacheBuffer;
  reg                 badvICacheBufferLock;
  wire                when_CSR_l173;
  wire                when_CSR_l176;
  reg        [4:0]    badvDCacheROBIdx;
  reg        [31:0]   badvDCacheBuffer;
  reg                 badvDCacheBufferLock;
  wire                when_CSR_l189;
  wire                when_CSR_l193;
  wire       [31:0]   _zz_io_interrupt_1;
  wire       [31:0]   _zz_io_swRead_value_113;
  wire       [31:0]   _zz_io_swRead_value_114;
  wire       [31:0]   _zz_io_swRead_value_115;
  wire       [31:0]   _zz_io_swRead_value_116;
  wire       [31:0]   _zz_io_swRead_value_117;
  wire       [31:0]   _zz_io_swRead_value_118;
  wire       [31:0]   _zz_io_swRead_value_119;
  wire       [31:0]   _zz_io_swRead_value_120;
  wire       [31:0]   _zz_io_swRead_value_121;
  wire       [31:0]   _zz_io_swRead_value_122;
  wire       [31:0]   _zz_io_swRead_value_123;
  wire       [30:0]   _zz_io_swRead_value_124;
  wire                when_CSR_l272;
  wire       [31:0]   _zz_io_swRead_value_125;
  wire       [31:0]   _zz_io_swRead_value_126;
  wire       [31:0]   _zz_io_swRead_value_127;
  wire                when_CSR_l289;
  wire                when_CSR_l303;
  wire                when_CSR_l305;
  wire                when_CSR_l313;
  wire                when_CSR_l314;
  function  zz_stableCounter_willIncrement(input dummy);
    begin
      zz_stableCounter_willIncrement = 1'b0;
      zz_stableCounter_willIncrement = 1'b1;
    end
  endfunction
  wire  _zz_1;

  assign _zz__zz_io_swRead_value_76 = 4'b1010;
  assign _zz_io_diffCSRBundle_ticlr = ticlr;
  assign _zz_stableCounter_valueNext_1 = stableCounter_willIncrement;
  assign _zz_stableCounter_valueNext = {63'd0, _zz_stableCounter_valueNext_1};
  assign _zz__zz_io_swRead_value_112 = (_zz_io_swRead_value_89 - _zz__zz_io_swRead_value_112_1);
  assign _zz__zz_io_swRead_value_112_2 = _zz_io_swRead_value_86;
  assign _zz__zz_io_swRead_value_112_1 = {31'd0, _zz__zz_io_swRead_value_112_2};
  assign _zz_intVec = {_zz_io_swRead_value_46,{_zz_io_swRead_value_45,{_zz_io_swRead_value_44,{_zz_io_swRead_value_43,{_zz_io_swRead_value_42,{_zz_io_swRead_value_41,{_zz_io_swRead_value_40,{_zz_io_swRead_value_39,_zz_io_swRead_value_38}}}}}}}};
  assign _zz_intVec_1 = {_zz_io_swRead_value_37,{_zz_io_swRead_value_36,{_zz_io_swRead_value_35,_zz_io_swRead_value_34}}};
  assign _zz__zz_io_interrupt_1 = {_zz_io_swRead_value_30,{_zz_io_swRead_value_29,{_zz_io_swRead_value_28,{_zz_io_swRead_value_27,{_zz_io_swRead_value_26,{_zz_io_interrupt,_zz_io_swRead_value_25}}}}}};
  assign _zz__zz_io_swRead_value_113 = {_zz_io_swRead_value_33,{_zz_io_swRead_value_32,_zz_io_swRead_value_31}};
  assign _zz__zz_io_swRead_value_114 = {_zz_io_swRead_value_37,{_zz_io_swRead_value_36,{_zz_io_swRead_value_35,_zz_io_swRead_value_34}}};
  assign _zz__zz_io_swRead_value_114_1 = {_zz_io_swRead_value_37,{_zz_io_swRead_value_36,{_zz_io_swRead_value_35,_zz_io_swRead_value_34}}};
  assign _zz__zz_io_swRead_value_115 = {_zz_io_swRead_value_46,{_zz_io_swRead_value_45,{_zz_io_swRead_value_44,{_zz_io_swRead_value_43,{_zz_io_swRead_value_42,{_zz_io_swRead_value_41,{_zz_io_swRead_value_40,{_zz_io_swRead_value_39,_zz_io_swRead_value_38}}}}}}}};
  assign _zz__zz_io_swRead_value_116 = {_zz_io_swRead_value_50,_zz_io_swRead_value_49};
  assign _zz__zz_io_swRead_value_117 = {_zz_io_swRead_value_55,{_zz_io_swRead_value_54,{_zz_io_swRead_value_53,{_zz_io_swRead_value_52,_zz_io_swRead_value_51}}}};
  assign _zz__zz_io_swRead_value_117_1 = {_zz_io_swRead_value_55,{_zz_io_swRead_value_54,{_zz_io_swRead_value_53,{_zz_io_swRead_value_52,_zz_io_swRead_value_51}}}};
  assign _zz__zz_io_swRead_value_118 = {_zz_io_swRead_value_57,_zz_io_swRead_value_56};
  assign _zz__zz_io_swRead_value_119 = {_zz_io_swRead_value_65,{_zz_io_swRead_value_64,{_zz_io_swRead_value_63,{_zz_io_swRead_value_62,{_zz_io_swRead_value_61,{_zz_io_swRead_value_60,{_zz_io_swRead_value_59,_zz_io_swRead_value_58}}}}}}};
  assign _zz__zz_io_swRead_value_119_1 = {_zz_io_swRead_value_65,{_zz_io_swRead_value_64,{_zz_io_swRead_value_63,{_zz_io_swRead_value_62,{_zz_io_swRead_value_61,{_zz_io_swRead_value_60,{_zz_io_swRead_value_59,_zz_io_swRead_value_58}}}}}}};
  assign _zz__zz_io_swRead_value_120 = {_zz_io_swRead_value_65,{_zz_io_swRead_value_64,{_zz_io_swRead_value_63,{_zz_io_swRead_value_62,{_zz_io_swRead_value_61,{_zz_io_swRead_value_60,{_zz_io_swRead_value_59,_zz_io_swRead_value_58}}}}}}};
  assign _zz__zz_io_swRead_value_120_1 = {_zz_io_swRead_value_65,{_zz_io_swRead_value_64,{_zz_io_swRead_value_63,{_zz_io_swRead_value_62,{_zz_io_swRead_value_61,{_zz_io_swRead_value_60,{_zz_io_swRead_value_59,_zz_io_swRead_value_58}}}}}}};
  assign _zz__zz_io_swRead_value_121 = {_zz_io_swRead_value_77,{_zz_io_swRead_value_76,{_zz_io_swRead_value_75,_zz_io_swRead_value_74}}};
  assign _zz__zz_io_swRead_value_122 = {_zz_io_swRead_value_79,_zz_io_swRead_value_78};
  assign _zz__zz_io_swRead_value_123 = {_zz_io_swRead_value_81,_zz_io_swRead_value_80};
  assign _zz__zz_io_swRead_value_124 = {_zz_io_swRead_value_93,{_zz_io_swRead_value_92,{_zz_io_swRead_value_91,_zz_io_swRead_value_90}}};
  assign _zz__zz_io_swRead_value_124_1 = {_zz_io_swRead_value_93,{_zz_io_swRead_value_92,{_zz_io_swRead_value_91,_zz_io_swRead_value_90}}};
  assign _zz__zz_io_swRead_value_125 = {_zz_io_swRead_value_95,_zz_io_swRead_value_94};
  assign _zz__zz_io_swRead_value_126 = {_zz_io_swRead_value_103,{_zz_io_swRead_value_102,{_zz_io_swRead_value_101,{_zz_io_swRead_value_100,{_zz_io_swRead_value_99,{_zz_io_swRead_value_98,{_zz_io_swRead_value_97,_zz_io_swRead_value_96}}}}}}};
  assign _zz__zz_io_swRead_value_126_1 = {_zz_io_swRead_value_103,{_zz_io_swRead_value_102,{_zz_io_swRead_value_101,{_zz_io_swRead_value_100,{_zz_io_swRead_value_99,{_zz_io_swRead_value_98,{_zz_io_swRead_value_97,_zz_io_swRead_value_96}}}}}}};
  assign _zz__zz_io_swRead_value_126_2 = {_zz_io_swRead_value_103,{_zz_io_swRead_value_102,{_zz_io_swRead_value_101,{_zz_io_swRead_value_100,{_zz_io_swRead_value_99,{_zz_io_swRead_value_98,{_zz_io_swRead_value_97,_zz_io_swRead_value_96}}}}}}};
  assign _zz__zz_io_swRead_value_127 = {_zz_io_swRead_value_111,{_zz_io_swRead_value_110,{_zz_io_swRead_value_109,{_zz_io_swRead_value_108,{_zz_io_swRead_value_107,{_zz_io_swRead_value_106,{_zz_io_swRead_value_105,_zz_io_swRead_value_104}}}}}}};
  assign _zz__zz_io_swRead_value_127_1 = {_zz_io_swRead_value_111,{_zz_io_swRead_value_110,{_zz_io_swRead_value_109,{_zz_io_swRead_value_108,{_zz_io_swRead_value_107,{_zz_io_swRead_value_106,{_zz_io_swRead_value_105,_zz_io_swRead_value_104}}}}}}};
  assign _zz__zz_io_swRead_value_127_2 = {_zz_io_swRead_value_111,{_zz_io_swRead_value_110,{_zz_io_swRead_value_109,{_zz_io_swRead_value_108,{_zz_io_swRead_value_107,{_zz_io_swRead_value_106,{_zz_io_swRead_value_105,_zz_io_swRead_value_104}}}}}}};
  assign _zz_when_CSR_l303_4 = 1'b1;
  assign _zz_when_CSR_l303_3 = {5'd0, _zz_when_CSR_l303_4};
  assign _zz_when_CSR_l303_7 = 2'b10;
  assign _zz_when_CSR_l303_6 = {4'd0, _zz_when_CSR_l303_7};
  assign _zz_when_CSR_l303_10 = 2'b11;
  assign _zz_when_CSR_l303_9 = {4'd0, _zz_when_CSR_l303_10};
  assign _zz_when_CSR_l303_12 = 3'b100;
  assign _zz_when_CSR_l303_11 = {3'd0, _zz_when_CSR_l303_12};
  assign _zz_when_CSR_l303_14 = 3'b111;
  assign _zz_when_CSR_l303_13 = {3'd0, _zz_when_CSR_l303_14};
  assign _zz_when_CSR_l313_1 = 4'b1000;
  assign _zz_when_CSR_l313 = {2'd0, _zz_when_CSR_l313_1};
  assign _zz_when_CSR_l313_3 = 4'b1001;
  assign _zz_when_CSR_l313_2 = {2'd0, _zz_when_CSR_l313_3};
  assign _zz_when_CSR_l303 = (io_ctrl_eCode == 6'h3f);
  assign _zz_when_CSR_l303_1 = (io_ctrl_eSubCode == 1'b0);
  assign _zz_when_CSR_l303_2 = (io_ctrl_eCode == _zz_when_CSR_l303_3);
  assign _zz_when_CSR_l303_5 = (io_ctrl_eSubCode == 1'b0);
  assign _zz_when_CSR_l303_8 = 1'b0;
  assign io_diffCSRBundle_crmd = {_zz_io_swRead_value_30,{_zz_io_swRead_value_29,{_zz_io_swRead_value_28,{_zz_io_swRead_value_27,{_zz_io_swRead_value_26,{_zz_io_interrupt,_zz_io_swRead_value_25}}}}}};
  assign io_diffCSRBundle_prmd = {_zz_io_swRead_value_33,{_zz_io_swRead_value_32,_zz_io_swRead_value_31}};
  assign io_diffCSRBundle_ecfg = {_zz_io_swRead_value_37,{_zz_io_swRead_value_36,{_zz_io_swRead_value_35,_zz_io_swRead_value_34}}};
  assign io_diffCSRBundle_estat = {_zz_io_swRead_value_46,{_zz_io_swRead_value_45,{_zz_io_swRead_value_44,{_zz_io_swRead_value_43,{_zz_io_swRead_value_42,{_zz_io_swRead_value_41,{_zz_io_swRead_value_40,{_zz_io_swRead_value_39,_zz_io_swRead_value_38}}}}}}}};
  assign io_diffCSRBundle_era = _zz_io_swRead_value_47;
  assign io_diffCSRBundle_badv = _zz_io_swRead_value_48;
  assign io_diffCSRBundle_eentry = {_zz_io_swRead_value_50,_zz_io_swRead_value_49};
  assign io_diffCSRBundle_tlbidx = {_zz_io_swRead_value_55,{_zz_io_swRead_value_54,{_zz_io_swRead_value_53,{_zz_io_swRead_value_52,_zz_io_swRead_value_51}}}};
  assign io_diffCSRBundle_tlbehi = {_zz_io_swRead_value_57,_zz_io_swRead_value_56};
  assign io_diffCSRBundle_tlbelo0 = {_zz_io_swRead_value_65,{_zz_io_swRead_value_64,{_zz_io_swRead_value_63,{_zz_io_swRead_value_62,{_zz_io_swRead_value_61,{_zz_io_swRead_value_60,{_zz_io_swRead_value_59,_zz_io_swRead_value_58}}}}}}};
  assign io_diffCSRBundle_tlbelo1 = {_zz_io_swRead_value_73,{_zz_io_swRead_value_72,{_zz_io_swRead_value_71,{_zz_io_swRead_value_70,{_zz_io_swRead_value_69,{_zz_io_swRead_value_68,{_zz_io_swRead_value_67,_zz_io_swRead_value_66}}}}}}};
  assign io_diffCSRBundle_asid = {_zz_io_swRead_value_77,{_zz_io_swRead_value_76,{_zz_io_swRead_value_75,_zz_io_swRead_value_74}}};
  assign io_diffCSRBundle_pgdl = {_zz_io_swRead_value_79,_zz_io_swRead_value_78};
  assign io_diffCSRBundle_pgdh = {_zz_io_swRead_value_81,_zz_io_swRead_value_80};
  assign io_diffCSRBundle_save0 = _zz_io_swRead_value_82;
  assign io_diffCSRBundle_save1 = _zz_io_swRead_value_83;
  assign io_diffCSRBundle_save2 = _zz_io_swRead_value_84;
  assign io_diffCSRBundle_save3 = _zz_io_swRead_value_85;
  assign io_diffCSRBundle_tid = _zz_io_counter_id;
  assign io_diffCSRBundle_tcfg = {_zz_io_swRead_value_88,{_zz_io_swRead_value_87,_zz_io_swRead_value_86}};
  assign io_diffCSRBundle_tval = _zz_io_swRead_value_89;
  assign io_diffCSRBundle_ticlr = {31'd0, _zz_io_diffCSRBundle_ticlr};
  assign io_diffCSRBundle_llbctl = {_zz_io_swRead_value_93,{_zz_io_swRead_value_92,{_zz_io_swRead_value_91,_zz_io_swRead_value_90}}};
  assign io_diffCSRBundle_tlbrentry = {_zz_io_swRead_value_95,_zz_io_swRead_value_94};
  assign io_diffCSRBundle_dmw0 = {_zz_io_swRead_value_103,{_zz_io_swRead_value_102,{_zz_io_swRead_value_101,{_zz_io_swRead_value_100,{_zz_io_swRead_value_99,{_zz_io_swRead_value_98,{_zz_io_swRead_value_97,_zz_io_swRead_value_96}}}}}}};
  assign io_diffCSRBundle_dmw1 = {_zz_io_swRead_value_111,{_zz_io_swRead_value_110,{_zz_io_swRead_value_109,{_zz_io_swRead_value_108,{_zz_io_swRead_value_107,{_zz_io_swRead_value_106,{_zz_io_swRead_value_105,_zz_io_swRead_value_104}}}}}}};
  assign _zz_1 = zz_stableCounter_willIncrement(1'b0);
  always @(*) stableCounter_willIncrement = _zz_1;
  assign stableCounter_willClear = 1'b0;
  assign stableCounter_willOverflowIfInc = (stableCounter_value == 64'hffffffffffffffff);
  assign stableCounter_willOverflow = (stableCounter_willOverflowIfInc && stableCounter_willIncrement);
  always @(*) begin
    stableCounter_valueNext = (stableCounter_value + _zz_stableCounter_valueNext);
    if(stableCounter_willClear) begin
      stableCounter_valueNext = 64'h0000000000000000;
    end
  end

  always @(*) begin
    ticlr = 1'b0;
    if(io_ctrl_writeCSR) begin
      case(csrWriteBuffer_address)
        14'h0044 : begin
          ticlr = csrWriteBuffer_value[0];
        end
        default : begin
        end
      endcase
    end
  end

  assign timeUp = ((_zz_io_swRead_value_89 == 32'h00000001) && _zz_io_swRead_value_86);
  assign when_CSR_l116 = (_zz_io_swRead_value_89 == 32'h00000000);
  assign when_CSR_l117 = (_zz_io_swRead_value_87 && _zz_io_swRead_value_86);
  always @(*) begin
    if(when_CSR_l116) begin
      if(when_CSR_l117) begin
        _zz_io_swRead_value_112 = {_zz_io_swRead_value_88,2'b00};
      end else begin
        _zz_io_swRead_value_112 = 32'h00000000;
      end
    end else begin
      _zz_io_swRead_value_112 = _zz__zz_io_swRead_value_112;
    end
  end

  assign intVec = (_zz_intVec[15 : 0] & _zz_intVec_1[15 : 0]);
  assign when_CSR_l139 = (io_swWrite_wen && (! csrWriteBufferLock));
  assign when_CSR_l143 = (io_swWrite_wen && (! io_flush));
  assign when_CSR_l156 = (io_llBitComm_wen && (! llbUpdateBufferLock));
  assign when_CSR_l159 = (io_llBitComm_wen && (! io_flush));
  assign when_CSR_l173 = (io_badvICache_wen && (! badvICacheBufferLock));
  assign when_CSR_l176 = (io_badvICache_wen && (! io_flush));
  assign when_CSR_l189 = (io_badvDCache_wen && (! badvDCacheBufferLock));
  assign when_CSR_l193 = (io_badvDCache_wen && (! io_flush));
  always @(*) begin
    case(io_swRead_address)
      14'h0000 : begin
        io_swRead_value = {_zz_io_swRead_value_30,{_zz_io_swRead_value_29,{_zz_io_swRead_value_28,{_zz_io_swRead_value_27,{_zz_io_swRead_value_26,{_zz_io_interrupt,_zz_io_swRead_value_25}}}}}};
      end
      14'h0001 : begin
        io_swRead_value = {_zz_io_swRead_value_33,{_zz_io_swRead_value_32,_zz_io_swRead_value_31}};
      end
      14'h0004 : begin
        io_swRead_value = {_zz_io_swRead_value_37,{_zz_io_swRead_value_36,{_zz_io_swRead_value_35,_zz_io_swRead_value_34}}};
      end
      14'h0005 : begin
        io_swRead_value = {_zz_io_swRead_value_46,{_zz_io_swRead_value_45,{_zz_io_swRead_value_44,{_zz_io_swRead_value_43,{_zz_io_swRead_value_42,{_zz_io_swRead_value_41,{_zz_io_swRead_value_40,{_zz_io_swRead_value_39,_zz_io_swRead_value_38}}}}}}}};
      end
      14'h0006 : begin
        io_swRead_value = _zz_io_swRead_value_47;
      end
      14'h0007 : begin
        io_swRead_value = _zz_io_swRead_value_48;
      end
      14'h000c : begin
        io_swRead_value = {_zz_io_swRead_value_50,_zz_io_swRead_value_49};
      end
      14'h0010 : begin
        io_swRead_value = {_zz_io_swRead_value_55,{_zz_io_swRead_value_54,{_zz_io_swRead_value_53,{_zz_io_swRead_value_52,_zz_io_swRead_value_51}}}};
      end
      14'h0011 : begin
        io_swRead_value = {_zz_io_swRead_value_57,_zz_io_swRead_value_56};
      end
      14'h0012 : begin
        io_swRead_value = {_zz_io_swRead_value_65,{_zz_io_swRead_value_64,{_zz_io_swRead_value_63,{_zz_io_swRead_value_62,{_zz_io_swRead_value_61,{_zz_io_swRead_value_60,{_zz_io_swRead_value_59,_zz_io_swRead_value_58}}}}}}};
      end
      14'h0013 : begin
        io_swRead_value = {_zz_io_swRead_value_73,{_zz_io_swRead_value_72,{_zz_io_swRead_value_71,{_zz_io_swRead_value_70,{_zz_io_swRead_value_69,{_zz_io_swRead_value_68,{_zz_io_swRead_value_67,_zz_io_swRead_value_66}}}}}}};
      end
      14'h0018 : begin
        io_swRead_value = {_zz_io_swRead_value_77,{_zz_io_swRead_value_76,{_zz_io_swRead_value_75,_zz_io_swRead_value_74}}};
      end
      14'h0019 : begin
        io_swRead_value = {_zz_io_swRead_value_79,_zz_io_swRead_value_78};
      end
      14'h001a : begin
        io_swRead_value = {_zz_io_swRead_value_81,_zz_io_swRead_value_80};
      end
      14'h001b : begin
        io_swRead_value = (_zz_io_swRead_value_48[31] ? {_zz_io_swRead_value_81,_zz_io_swRead_value_80} : {_zz_io_swRead_value_79,_zz_io_swRead_value_78});
      end
      14'h0020 : begin
        io_swRead_value = 32'h00000000;
      end
      14'h0030 : begin
        io_swRead_value = _zz_io_swRead_value_82;
      end
      14'h0031 : begin
        io_swRead_value = _zz_io_swRead_value_83;
      end
      14'h0032 : begin
        io_swRead_value = _zz_io_swRead_value_84;
      end
      14'h0033 : begin
        io_swRead_value = _zz_io_swRead_value_85;
      end
      14'h0040 : begin
        io_swRead_value = _zz_io_counter_id;
      end
      14'h0041 : begin
        io_swRead_value = {_zz_io_swRead_value_88,{_zz_io_swRead_value_87,_zz_io_swRead_value_86}};
      end
      14'h0042 : begin
        io_swRead_value = _zz_io_swRead_value_89;
      end
      14'h0044 : begin
        io_swRead_value = 32'h00000000;
      end
      14'h0060 : begin
        io_swRead_value = {_zz_io_swRead_value_93,{_zz_io_swRead_value_92,{_zz_io_swRead_value_91,_zz_io_swRead_value_90}}};
      end
      14'h0088 : begin
        io_swRead_value = {_zz_io_swRead_value_95,_zz_io_swRead_value_94};
      end
      14'h0180 : begin
        io_swRead_value = {_zz_io_swRead_value_103,{_zz_io_swRead_value_102,{_zz_io_swRead_value_101,{_zz_io_swRead_value_100,{_zz_io_swRead_value_99,{_zz_io_swRead_value_98,{_zz_io_swRead_value_97,_zz_io_swRead_value_96}}}}}}};
      end
      14'h0181 : begin
        io_swRead_value = {_zz_io_swRead_value_111,{_zz_io_swRead_value_110,{_zz_io_swRead_value_109,{_zz_io_swRead_value_108,{_zz_io_swRead_value_107,{_zz_io_swRead_value_106,{_zz_io_swRead_value_105,_zz_io_swRead_value_104}}}}}}};
      end
      default : begin
        io_swRead_value = 32'h00000000;
      end
    endcase
  end

  assign _zz_io_interrupt_1 = {_zz__zz_io_interrupt_1[31 : 9],csrWriteBuffer_value[8 : 0]};
  assign _zz_io_swRead_value_113 = {_zz__zz_io_swRead_value_113[31 : 3],csrWriteBuffer_value[2 : 0]};
  assign _zz_io_swRead_value_114 = {{{_zz__zz_io_swRead_value_114[31 : 13],csrWriteBuffer_value[12 : 11]},_zz__zz_io_swRead_value_114_1[10]},csrWriteBuffer_value[9 : 0]};
  assign _zz_io_swRead_value_115 = {_zz__zz_io_swRead_value_115[31 : 2],csrWriteBuffer_value[1 : 0]};
  assign _zz_io_swRead_value_116 = {csrWriteBuffer_value[31 : 6],_zz__zz_io_swRead_value_116[5 : 0]};
  assign _zz_io_swRead_value_117 = {{{{csrWriteBuffer_value[31],_zz__zz_io_swRead_value_117[30]},csrWriteBuffer_value[29 : 24]},_zz__zz_io_swRead_value_117_1[23 : 2]},csrWriteBuffer_value[1 : 0]};
  assign _zz_io_swRead_value_118 = {csrWriteBuffer_value[31 : 13],_zz__zz_io_swRead_value_118[12 : 0]};
  assign _zz_io_swRead_value_119 = {{{_zz__zz_io_swRead_value_119[31 : 28],csrWriteBuffer_value[27 : 8]},_zz__zz_io_swRead_value_119_1[7]},csrWriteBuffer_value[6 : 0]};
  assign _zz_io_swRead_value_120 = {{{_zz__zz_io_swRead_value_120[31 : 28],csrWriteBuffer_value[27 : 8]},_zz__zz_io_swRead_value_120_1[7]},csrWriteBuffer_value[6 : 0]};
  assign _zz_io_swRead_value_121 = {_zz__zz_io_swRead_value_121[31 : 10],csrWriteBuffer_value[9 : 0]};
  assign _zz_io_swRead_value_122 = {csrWriteBuffer_value[31 : 12],_zz__zz_io_swRead_value_122[11 : 0]};
  assign _zz_io_swRead_value_123 = {csrWriteBuffer_value[31 : 12],_zz__zz_io_swRead_value_123[11 : 0]};
  assign _zz_io_swRead_value_124 = {{_zz__zz_io_swRead_value_124[31 : 3],csrWriteBuffer_value[2]},_zz__zz_io_swRead_value_124_1[1]};
  assign when_CSR_l272 = csrWriteBuffer_value[1];
  assign _zz_io_swRead_value_125 = {csrWriteBuffer_value[31 : 6],_zz__zz_io_swRead_value_125[5 : 0]};
  assign _zz_io_swRead_value_126 = {{{{{{csrWriteBuffer_value[31 : 29],_zz__zz_io_swRead_value_126[28]},csrWriteBuffer_value[27 : 25]},_zz__zz_io_swRead_value_126_1[24 : 6]},csrWriteBuffer_value[5 : 3]},_zz__zz_io_swRead_value_126_2[2 : 1]},csrWriteBuffer_value[0]};
  assign _zz_io_swRead_value_127 = {{{{{{csrWriteBuffer_value[31 : 29],_zz__zz_io_swRead_value_127[28]},csrWriteBuffer_value[27 : 25]},_zz__zz_io_swRead_value_127_1[24 : 6]},csrWriteBuffer_value[5 : 3]},_zz__zz_io_swRead_value_127_2[2 : 1]},csrWriteBuffer_value[0]};
  assign when_CSR_l289 = (io_ctrl_normalException || io_ctrl_tlbrException);
  assign when_CSR_l303 = ((((((_zz_when_CSR_l303 && _zz_when_CSR_l303_1) || (_zz_when_CSR_l303_2 && _zz_when_CSR_l303_5)) || ((io_ctrl_eCode == _zz_when_CSR_l303_6) && (io_ctrl_eSubCode == _zz_when_CSR_l303_8))) || ((io_ctrl_eCode == _zz_when_CSR_l303_9) && (io_ctrl_eSubCode == 1'b0))) || ((io_ctrl_eCode == _zz_when_CSR_l303_11) && (io_ctrl_eSubCode == 1'b0))) || ((io_ctrl_eCode == _zz_when_CSR_l303_13) && (io_ctrl_eSubCode == 1'b0)));
  assign when_CSR_l305 = ((io_ctrl_eROBIdx == badvDCacheROBIdx) && badvDCacheBufferLock);
  assign when_CSR_l313 = (((io_ctrl_eCode == _zz_when_CSR_l313) && (io_ctrl_eSubCode == 1'b0)) || ((io_ctrl_eCode == _zz_when_CSR_l313_2) && (io_ctrl_eSubCode == 1'b0)));
  assign when_CSR_l314 = ((io_ctrl_eROBIdx == badvDCacheROBIdx) && badvDCacheBufferLock);
  assign io_interrupt = (_zz_io_interrupt && (|intVec));
  assign _zz_when_Cache_l83 = _zz_io_swRead_value_25;
  assign io_counter_id = _zz_io_counter_id;
  assign io_counter_value = stableCounter_value;
  assign io_llBitComm_actualAddr = llAddr;
  assign _zz_scMatchHit = _zz_io_swRead_value_90;
  assign io_tlbCSRInfo_asid = _zz_io_swRead_value_74;
  assign _zz_io_iCacheReq_pageInfo_plv = _zz_io_swRead_value_25;
  assign _zz_when_TLB_l177 = _zz_io_swRead_value_26;
  assign _zz_when_TLB_l177_1 = _zz_io_swRead_value_27;
  assign _zz_io_iCacheReq_pageInfo_mat = _zz_io_swRead_value_28;
  assign _zz_io_dCacheReq_pageInfo_mat = _zz_io_swRead_value_29;
  assign _zz_when_TLB_l178 = _zz_io_swRead_value_96;
  assign _zz_when_TLB_l178_1 = _zz_io_swRead_value_98;
  assign _zz_io_iCacheReq_pageInfo_mat_1 = _zz_io_swRead_value_99;
  assign _zz_io_iCacheReq_pageInfo_ppn = _zz_io_swRead_value_101;
  assign _zz_when_TLB_l178_2 = _zz_io_swRead_value_103;
  assign _zz_when_TLB_l185 = _zz_io_swRead_value_104;
  assign _zz_when_TLB_l185_1 = _zz_io_swRead_value_106;
  assign _zz_io_iCacheReq_pageInfo_mat_2 = _zz_io_swRead_value_107;
  assign _zz_io_iCacheReq_pageInfo_ppn_1 = _zz_io_swRead_value_109;
  assign _zz_when_TLB_l185_2 = _zz_io_swRead_value_111;
  assign _zz_entryToFill_e = _zz_io_swRead_value_44;
  assign _zz_io_csrWrite_asid = _zz_io_swRead_value_51;
  assign _zz_io_swRead_value = _zz_io_swRead_value_52;
  assign _zz_entryToFill_ps = _zz_io_swRead_value_53;
  assign _zz_io_swRead_value_1 = _zz_io_swRead_value_54;
  assign _zz_entryToFill_e_1 = _zz_io_swRead_value_55;
  assign _zz_entryToFill_vppn = _zz_io_swRead_value_57;
  assign _zz_entryToFill_pp0_v = _zz_io_swRead_value_58;
  assign _zz_entryToFill_pp0_d = _zz_io_swRead_value_59;
  assign _zz_entryToFill_pp0_plv = _zz_io_swRead_value_60;
  assign _zz_entryToFill_pp0_mat = _zz_io_swRead_value_61;
  assign _zz_entryToFill_g = _zz_io_swRead_value_62;
  assign _zz_entryToFill_pp0_ppn = _zz_io_swRead_value_64;
  assign _zz_entryToFill_pp1_v = _zz_io_swRead_value_66;
  assign _zz_entryToFill_pp1_d = _zz_io_swRead_value_67;
  assign _zz_entryToFill_pp1_plv = _zz_io_swRead_value_68;
  assign _zz_entryToFill_pp1_mat = _zz_io_swRead_value_69;
  assign _zz_entryToFill_g_1 = _zz_io_swRead_value_70;
  assign _zz_entryToFill_pp1_ppn = _zz_io_swRead_value_72;
  assign io_ctrl_era = _zz_io_swRead_value_47;
  assign io_ctrl_eentry = {_zz_io_swRead_value_50,_zz_io_swRead_value_49};
  assign io_ctrl_tlbrentry = {_zz_io_swRead_value_95,_zz_io_swRead_value_94};
  always @(posedge aclk) begin
    if(!aresetn) begin
      _zz_io_swRead_value_25 <= 2'b00;
      _zz_io_interrupt <= 1'b0;
      _zz_io_swRead_value_26 <= 1'b1;
      _zz_io_swRead_value_27 <= 1'b0;
      _zz_io_swRead_value_28 <= 2'b00;
      _zz_io_swRead_value_29 <= 2'b00;
      _zz_io_swRead_value_30 <= 23'h000000;
      _zz_io_swRead_value_31 <= 2'b00;
      _zz_io_swRead_value_32 <= 1'b0;
      _zz_io_swRead_value_33 <= 29'h00000000;
      _zz_io_swRead_value_34 <= 10'h000;
      _zz_io_swRead_value_35 <= 1'b0;
      _zz_io_swRead_value_36 <= 2'b00;
      _zz_io_swRead_value_37 <= 19'h00000;
      _zz_io_swRead_value_38 <= 2'b00;
      _zz_io_swRead_value_39 <= 8'h00;
      _zz_io_swRead_value_40 <= 1'b0;
      _zz_io_swRead_value_41 <= 1'b0;
      _zz_io_swRead_value_42 <= 1'b0;
      _zz_io_swRead_value_43 <= 3'b000;
      _zz_io_swRead_value_44 <= 6'h00;
      _zz_io_swRead_value_45 <= 9'h000;
      _zz_io_swRead_value_46 <= 1'b0;
      _zz_io_swRead_value_47 <= 32'h00000000;
      _zz_io_swRead_value_48 <= 32'h00000000;
      _zz_io_swRead_value_49 <= 6'h00;
      _zz_io_swRead_value_50 <= 26'h0000000;
      _zz_io_swRead_value_51 <= 2'b00;
      _zz_io_swRead_value_52 <= 22'h000000;
      _zz_io_swRead_value_53 <= 6'h00;
      _zz_io_swRead_value_54 <= 1'b0;
      _zz_io_swRead_value_55 <= 1'b0;
      _zz_io_swRead_value_56 <= 13'h0000;
      _zz_io_swRead_value_57 <= 19'h00000;
      _zz_io_swRead_value_58 <= 1'b0;
      _zz_io_swRead_value_59 <= 1'b0;
      _zz_io_swRead_value_60 <= 2'b00;
      _zz_io_swRead_value_61 <= 2'b00;
      _zz_io_swRead_value_62 <= 1'b0;
      _zz_io_swRead_value_63 <= 1'b0;
      _zz_io_swRead_value_64 <= 20'h00000;
      _zz_io_swRead_value_65 <= 4'b0000;
      _zz_io_swRead_value_66 <= 1'b0;
      _zz_io_swRead_value_67 <= 1'b0;
      _zz_io_swRead_value_68 <= 2'b00;
      _zz_io_swRead_value_69 <= 2'b00;
      _zz_io_swRead_value_70 <= 1'b0;
      _zz_io_swRead_value_71 <= 1'b0;
      _zz_io_swRead_value_72 <= 20'h00000;
      _zz_io_swRead_value_73 <= 4'b0000;
      _zz_io_swRead_value_74 <= 10'h000;
      _zz_io_swRead_value_75 <= 6'h00;
      _zz_io_swRead_value_76 <= {4'd0, _zz__zz_io_swRead_value_76};
      _zz_io_swRead_value_77 <= 8'h00;
      _zz_io_swRead_value_78 <= 12'h000;
      _zz_io_swRead_value_79 <= 20'h00000;
      _zz_io_swRead_value_80 <= 12'h000;
      _zz_io_swRead_value_81 <= 20'h00000;
      _zz_io_swRead_value_82 <= 32'h00000000;
      _zz_io_swRead_value_83 <= 32'h00000000;
      _zz_io_swRead_value_84 <= 32'h00000000;
      _zz_io_swRead_value_85 <= 32'h00000000;
      _zz_io_counter_id <= 32'h00000000;
      _zz_io_swRead_value_86 <= 1'b0;
      _zz_io_swRead_value_87 <= 1'b0;
      _zz_io_swRead_value_88 <= 30'h00000000;
      _zz_io_swRead_value_89 <= {30'h00000000,2'b00};
      _zz_io_swRead_value_90 <= 1'b0;
      _zz_io_swRead_value_91 <= 1'b0;
      _zz_io_swRead_value_92 <= 1'b0;
      _zz_io_swRead_value_93 <= 29'h00000000;
      _zz_io_swRead_value_94 <= 6'h00;
      _zz_io_swRead_value_95 <= 26'h0000000;
      _zz_io_swRead_value_96 <= 1'b0;
      _zz_io_swRead_value_97 <= 2'b00;
      _zz_io_swRead_value_98 <= 1'b0;
      _zz_io_swRead_value_99 <= 2'b00;
      _zz_io_swRead_value_100 <= 19'h00000;
      _zz_io_swRead_value_101 <= 3'b000;
      _zz_io_swRead_value_102 <= 1'b0;
      _zz_io_swRead_value_103 <= 3'b000;
      _zz_io_swRead_value_104 <= 1'b0;
      _zz_io_swRead_value_105 <= 2'b00;
      _zz_io_swRead_value_106 <= 1'b0;
      _zz_io_swRead_value_107 <= 2'b00;
      _zz_io_swRead_value_108 <= 19'h00000;
      _zz_io_swRead_value_109 <= 3'b000;
      _zz_io_swRead_value_110 <= 1'b0;
      _zz_io_swRead_value_111 <= 3'b000;
      stableCounter_value <= 64'h0000000000000000;
      csrWriteBuffer_value <= 32'h00000000;
      csrWriteBuffer_address <= 14'h0000;
      csrWriteBufferLock <= 1'b0;
      llAddr <= 32'h00000000;
      llbUpdateBuffer <= 32'h00000000;
      llbUpdateBufferLock <= 1'b0;
      badvICacheBuffer <= 32'h00000000;
      badvICacheBufferLock <= 1'b0;
      badvDCacheROBIdx <= 5'h00;
      badvDCacheBuffer <= 32'h00000000;
      badvDCacheBufferLock <= 1'b0;
    end else begin
      stableCounter_value <= stableCounter_valueNext;
      _zz_io_swRead_value_89 <= _zz_io_swRead_value_112;
      _zz_io_swRead_value_39 <= io_extInt;
      _zz_io_swRead_value_41 <= ((timeUp || _zz_io_swRead_value_41) && (! ticlr));
      if(when_CSR_l139) begin
        csrWriteBuffer_value <= io_swWrite_value;
        csrWriteBuffer_address <= io_swWrite_address;
      end
      if(when_CSR_l143) begin
        csrWriteBufferLock <= 1'b1;
      end
      if(io_flush) begin
        csrWriteBufferLock <= 1'b0;
      end
      if(when_CSR_l156) begin
        llbUpdateBuffer <= io_llBitComm_toUpdateAddr;
      end
      if(when_CSR_l159) begin
        llbUpdateBufferLock <= 1'b1;
      end
      if(io_flush) begin
        llbUpdateBufferLock <= 1'b0;
      end
      if(io_ctrl_llBitUpdate) begin
        llAddr <= llbUpdateBuffer;
      end
      if(when_CSR_l173) begin
        badvICacheBuffer <= io_badvICache_vaddr;
      end
      if(when_CSR_l176) begin
        badvICacheBufferLock <= 1'b1;
      end
      if(io_flush) begin
        badvICacheBufferLock <= 1'b0;
      end
      if(when_CSR_l189) begin
        badvDCacheROBIdx <= io_badvDCache_robIdx;
        badvDCacheBuffer <= io_badvDCache_vaddr;
      end
      if(when_CSR_l193) begin
        badvDCacheBufferLock <= 1'b1;
      end
      if(io_flush) begin
        badvDCacheBufferLock <= 1'b0;
      end
      if(io_ctrl_writeCSR) begin
        case(csrWriteBuffer_address)
          14'h0000 : begin
            _zz_io_swRead_value_25 <= _zz_io_interrupt_1[1 : 0];
            _zz_io_interrupt <= _zz_io_interrupt_1[2];
            _zz_io_swRead_value_26 <= _zz_io_interrupt_1[3];
            _zz_io_swRead_value_27 <= _zz_io_interrupt_1[4];
            _zz_io_swRead_value_28 <= _zz_io_interrupt_1[6 : 5];
            _zz_io_swRead_value_29 <= _zz_io_interrupt_1[8 : 7];
            _zz_io_swRead_value_30 <= _zz_io_interrupt_1[31 : 9];
          end
          14'h0001 : begin
            _zz_io_swRead_value_31 <= _zz_io_swRead_value_113[1 : 0];
            _zz_io_swRead_value_32 <= _zz_io_swRead_value_113[2];
            _zz_io_swRead_value_33 <= _zz_io_swRead_value_113[31 : 3];
          end
          14'h0004 : begin
            _zz_io_swRead_value_34 <= _zz_io_swRead_value_114[9 : 0];
            _zz_io_swRead_value_35 <= _zz_io_swRead_value_114[10];
            _zz_io_swRead_value_36 <= _zz_io_swRead_value_114[12 : 11];
            _zz_io_swRead_value_37 <= _zz_io_swRead_value_114[31 : 13];
          end
          14'h0005 : begin
            _zz_io_swRead_value_38 <= _zz_io_swRead_value_115[1 : 0];
            _zz_io_swRead_value_39 <= _zz_io_swRead_value_115[9 : 2];
            _zz_io_swRead_value_40 <= _zz_io_swRead_value_115[10];
            _zz_io_swRead_value_41 <= _zz_io_swRead_value_115[11];
            _zz_io_swRead_value_42 <= _zz_io_swRead_value_115[12];
            _zz_io_swRead_value_43 <= _zz_io_swRead_value_115[15 : 13];
            _zz_io_swRead_value_44 <= _zz_io_swRead_value_115[21 : 16];
            _zz_io_swRead_value_45 <= _zz_io_swRead_value_115[30 : 22];
            _zz_io_swRead_value_46 <= _zz_io_swRead_value_115[31];
          end
          14'h0006 : begin
            _zz_io_swRead_value_47 <= csrWriteBuffer_value[31 : 0];
          end
          14'h0007 : begin
            _zz_io_swRead_value_48 <= csrWriteBuffer_value[31 : 0];
          end
          14'h000c : begin
            _zz_io_swRead_value_49 <= _zz_io_swRead_value_116[5 : 0];
            _zz_io_swRead_value_50 <= _zz_io_swRead_value_116[31 : 6];
          end
          14'h0010 : begin
            _zz_io_swRead_value_51 <= _zz_io_swRead_value_117[1 : 0];
            _zz_io_swRead_value_52 <= _zz_io_swRead_value_117[23 : 2];
            _zz_io_swRead_value_53 <= _zz_io_swRead_value_117[29 : 24];
            _zz_io_swRead_value_54 <= _zz_io_swRead_value_117[30];
            _zz_io_swRead_value_55 <= _zz_io_swRead_value_117[31];
          end
          14'h0011 : begin
            _zz_io_swRead_value_56 <= _zz_io_swRead_value_118[12 : 0];
            _zz_io_swRead_value_57 <= _zz_io_swRead_value_118[31 : 13];
          end
          14'h0012 : begin
            _zz_io_swRead_value_58 <= _zz_io_swRead_value_119[0];
            _zz_io_swRead_value_59 <= _zz_io_swRead_value_119[1];
            _zz_io_swRead_value_60 <= _zz_io_swRead_value_119[3 : 2];
            _zz_io_swRead_value_61 <= _zz_io_swRead_value_119[5 : 4];
            _zz_io_swRead_value_62 <= _zz_io_swRead_value_119[6];
            _zz_io_swRead_value_63 <= _zz_io_swRead_value_119[7];
            _zz_io_swRead_value_64 <= _zz_io_swRead_value_119[27 : 8];
            _zz_io_swRead_value_65 <= _zz_io_swRead_value_119[31 : 28];
          end
          14'h0013 : begin
            _zz_io_swRead_value_66 <= _zz_io_swRead_value_120[0];
            _zz_io_swRead_value_67 <= _zz_io_swRead_value_120[1];
            _zz_io_swRead_value_68 <= _zz_io_swRead_value_120[3 : 2];
            _zz_io_swRead_value_69 <= _zz_io_swRead_value_120[5 : 4];
            _zz_io_swRead_value_70 <= _zz_io_swRead_value_120[6];
            _zz_io_swRead_value_71 <= _zz_io_swRead_value_120[7];
            _zz_io_swRead_value_72 <= _zz_io_swRead_value_120[27 : 8];
            _zz_io_swRead_value_73 <= _zz_io_swRead_value_120[31 : 28];
          end
          14'h0018 : begin
            _zz_io_swRead_value_74 <= _zz_io_swRead_value_121[9 : 0];
            _zz_io_swRead_value_75 <= _zz_io_swRead_value_121[15 : 10];
            _zz_io_swRead_value_76 <= _zz_io_swRead_value_121[23 : 16];
            _zz_io_swRead_value_77 <= _zz_io_swRead_value_121[31 : 24];
          end
          14'h0019 : begin
            _zz_io_swRead_value_78 <= _zz_io_swRead_value_122[11 : 0];
            _zz_io_swRead_value_79 <= _zz_io_swRead_value_122[31 : 12];
          end
          14'h001a : begin
            _zz_io_swRead_value_80 <= _zz_io_swRead_value_123[11 : 0];
            _zz_io_swRead_value_81 <= _zz_io_swRead_value_123[31 : 12];
          end
          14'h0030 : begin
            _zz_io_swRead_value_82 <= csrWriteBuffer_value[31 : 0];
          end
          14'h0031 : begin
            _zz_io_swRead_value_83 <= csrWriteBuffer_value[31 : 0];
          end
          14'h0032 : begin
            _zz_io_swRead_value_84 <= csrWriteBuffer_value[31 : 0];
          end
          14'h0033 : begin
            _zz_io_swRead_value_85 <= csrWriteBuffer_value[31 : 0];
          end
          14'h0040 : begin
            _zz_io_counter_id <= csrWriteBuffer_value[31 : 0];
          end
          14'h0041 : begin
            _zz_io_swRead_value_86 <= csrWriteBuffer_value[0];
            _zz_io_swRead_value_87 <= csrWriteBuffer_value[1];
            _zz_io_swRead_value_88 <= csrWriteBuffer_value[31 : 2];
          end
          14'h0060 : begin
            _zz_io_swRead_value_91 <= _zz_io_swRead_value_124[0];
            _zz_io_swRead_value_92 <= _zz_io_swRead_value_124[1];
            _zz_io_swRead_value_93[28 : 0] <= _zz_io_swRead_value_124[30 : 2];
            if(when_CSR_l272) begin
              _zz_io_swRead_value_90 <= 1'b0;
            end
          end
          14'h0088 : begin
            _zz_io_swRead_value_94 <= _zz_io_swRead_value_125[5 : 0];
            _zz_io_swRead_value_95 <= _zz_io_swRead_value_125[31 : 6];
          end
          14'h0180 : begin
            _zz_io_swRead_value_96 <= _zz_io_swRead_value_126[0];
            _zz_io_swRead_value_97 <= _zz_io_swRead_value_126[2 : 1];
            _zz_io_swRead_value_98 <= _zz_io_swRead_value_126[3];
            _zz_io_swRead_value_99 <= _zz_io_swRead_value_126[5 : 4];
            _zz_io_swRead_value_100 <= _zz_io_swRead_value_126[24 : 6];
            _zz_io_swRead_value_101 <= _zz_io_swRead_value_126[27 : 25];
            _zz_io_swRead_value_102 <= _zz_io_swRead_value_126[28];
            _zz_io_swRead_value_103 <= _zz_io_swRead_value_126[31 : 29];
          end
          14'h0181 : begin
            _zz_io_swRead_value_104 <= _zz_io_swRead_value_127[0];
            _zz_io_swRead_value_105 <= _zz_io_swRead_value_127[2 : 1];
            _zz_io_swRead_value_106 <= _zz_io_swRead_value_127[3];
            _zz_io_swRead_value_107 <= _zz_io_swRead_value_127[5 : 4];
            _zz_io_swRead_value_108 <= _zz_io_swRead_value_127[24 : 6];
            _zz_io_swRead_value_109 <= _zz_io_swRead_value_127[27 : 25];
            _zz_io_swRead_value_110 <= _zz_io_swRead_value_127[28];
            _zz_io_swRead_value_111 <= _zz_io_swRead_value_127[31 : 29];
          end
          default : begin
          end
        endcase
      end
      if(io_ctrl_ertn) begin
        _zz_io_swRead_value_25 <= _zz_io_swRead_value_31;
        _zz_io_interrupt <= _zz_io_swRead_value_32;
        _zz_io_swRead_value_26 <= ((_zz_io_swRead_value_44 == 6'h3f) ? 1'b0 : _zz_io_swRead_value_26);
        _zz_io_swRead_value_27 <= ((_zz_io_swRead_value_44 == 6'h3f) ? 1'b1 : _zz_io_swRead_value_27);
        _zz_io_swRead_value_90 <= (_zz_io_swRead_value_92 ? _zz_io_swRead_value_90 : 1'b0);
        _zz_io_swRead_value_92 <= 1'b0;
      end
      if(when_CSR_l289) begin
        _zz_io_swRead_value_31 <= _zz_io_swRead_value_25;
        _zz_io_swRead_value_32 <= _zz_io_interrupt;
        _zz_io_swRead_value_25 <= 2'b00;
        _zz_io_interrupt <= 1'b0;
        _zz_io_swRead_value_47 <= io_ctrl_epc;
        _zz_io_swRead_value_44 <= io_ctrl_eCode;
        _zz_io_swRead_value_45 <= {8'd0, io_ctrl_eSubCode};
        if(when_CSR_l303) begin
          if(when_CSR_l305) begin
            _zz_io_swRead_value_48 <= badvDCacheBuffer;
            _zz_io_swRead_value_57 <= badvDCacheBuffer[31 : 13];
          end else begin
            _zz_io_swRead_value_48 <= badvICacheBuffer;
          end
        end
        if(when_CSR_l313) begin
          if(when_CSR_l314) begin
            _zz_io_swRead_value_48 <= badvDCacheBuffer;
          end else begin
            _zz_io_swRead_value_48 <= badvICacheBuffer;
          end
        end
        if(io_ctrl_tlbrException) begin
          _zz_io_swRead_value_26 <= 1'b1;
          _zz_io_swRead_value_27 <= 1'b0;
        end
      end
      if(io_tlbCSRWrite_idxWen) begin
        _zz_io_swRead_value_51 <= _zz_io_swRead_value_2;
        _zz_io_swRead_value_52 <= _zz_io_swRead_value_3;
        _zz_io_swRead_value_53 <= _zz_io_swRead_value_4;
        _zz_io_swRead_value_54 <= _zz_io_swRead_value_5;
        _zz_io_swRead_value_55 <= _zz_io_swRead_value_6;
      end
      if(io_tlbCSRWrite_entryWen) begin
        _zz_io_swRead_value_56 <= _zz_io_swRead_value_7;
        _zz_io_swRead_value_57 <= _zz_io_swRead_value_8;
        _zz_io_swRead_value_58 <= _zz_io_swRead_value_9;
        _zz_io_swRead_value_59 <= _zz_io_swRead_value_10;
        _zz_io_swRead_value_60 <= _zz_io_swRead_value_11;
        _zz_io_swRead_value_61 <= _zz_io_swRead_value_12;
        _zz_io_swRead_value_62 <= _zz_io_swRead_value_13;
        _zz_io_swRead_value_63 <= _zz_io_swRead_value_14;
        _zz_io_swRead_value_64 <= _zz_io_swRead_value_15;
        _zz_io_swRead_value_65 <= _zz_io_swRead_value_16;
        _zz_io_swRead_value_66 <= _zz_io_swRead_value_17;
        _zz_io_swRead_value_67 <= _zz_io_swRead_value_18;
        _zz_io_swRead_value_68 <= _zz_io_swRead_value_19;
        _zz_io_swRead_value_69 <= _zz_io_swRead_value_20;
        _zz_io_swRead_value_70 <= _zz_io_swRead_value_21;
        _zz_io_swRead_value_71 <= _zz_io_swRead_value_22;
        _zz_io_swRead_value_72 <= _zz_io_swRead_value_23;
        _zz_io_swRead_value_73 <= _zz_io_swRead_value_24;
        _zz_io_swRead_value_74 <= io_tlbCSRWrite_asid;
      end
    end
  end


endmodule

module ROB (
  input  wire [1:0]    io_dispatch_allowMask,
  output wire [1:0]    io_dispatch_availMask,
  output wire [4:0]    io_dispatch_robIdx_0,
  output wire [4:0]    io_dispatch_robIdx_1,
  input  wire [31:0]   io_dispatch_pc_0,
  input  wire [31:0]   io_dispatch_pc_1,
  input  wire [4:0]    io_dispatch_ard_0,
  input  wire [4:0]    io_dispatch_ard_1,
  input  wire [5:0]    io_dispatch_prd_0,
  input  wire [5:0]    io_dispatch_prd_1,
  input  wire [5:0]    io_dispatch_pprd_0,
  input  wire [5:0]    io_dispatch_pprd_1,
  input  wire [3:0]    io_dispatch_specialOp_0,
  input  wire [3:0]    io_dispatch_specialOp_1,
  input  wire [4:0]    io_commit_0_robIdx,
  input  wire [31:0]   io_commit_0_branchResult_targetPC,
  input  wire          io_commit_0_branchResult_branchResult,
  input  wire          io_commit_0_branchResult_predictFail,
  input  wire          io_commit_0_exceptionInfo_exception,
  input  wire [5:0]    io_commit_0_exceptionInfo_eCode,
  input  wire [0:0]    io_commit_0_exceptionInfo_eSubCode,
  input  wire          io_commit_0_valid,
  input  wire [4:0]    io_commit_1_robIdx,
  input  wire [31:0]   io_commit_1_branchResult_targetPC,
  input  wire          io_commit_1_branchResult_branchResult,
  input  wire          io_commit_1_branchResult_predictFail,
  input  wire          io_commit_1_exceptionInfo_exception,
  input  wire [5:0]    io_commit_1_exceptionInfo_eCode,
  input  wire [0:0]    io_commit_1_exceptionInfo_eSubCode,
  input  wire          io_commit_1_valid,
  input  wire [4:0]    io_commit_2_robIdx,
  input  wire [31:0]   io_commit_2_branchResult_targetPC,
  input  wire          io_commit_2_branchResult_branchResult,
  input  wire          io_commit_2_branchResult_predictFail,
  input  wire          io_commit_2_exceptionInfo_exception,
  input  wire [5:0]    io_commit_2_exceptionInfo_eCode,
  input  wire [0:0]    io_commit_2_exceptionInfo_eSubCode,
  input  wire          io_commit_2_valid,
  input  wire [4:0]    io_commit_3_robIdx,
  input  wire [31:0]   io_commit_3_branchResult_targetPC,
  input  wire          io_commit_3_branchResult_branchResult,
  input  wire          io_commit_3_branchResult_predictFail,
  input  wire          io_commit_3_exceptionInfo_exception,
  input  wire [5:0]    io_commit_3_exceptionInfo_eCode,
  input  wire [0:0]    io_commit_3_exceptionInfo_eSubCode,
  input  wire          io_commit_3_valid,
  input  wire [4:0]    io_commit_4_robIdx,
  input  wire [31:0]   io_commit_4_branchResult_targetPC,
  input  wire          io_commit_4_branchResult_branchResult,
  input  wire          io_commit_4_branchResult_predictFail,
  input  wire          io_commit_4_exceptionInfo_exception,
  input  wire [5:0]    io_commit_4_exceptionInfo_eCode,
  input  wire [0:0]    io_commit_4_exceptionInfo_eSubCode,
  input  wire          io_commit_4_valid,
  output wire [4:0]    io_retireARAT_0_ard,
  output wire [5:0]    io_retireARAT_0_prd,
  output wire          io_retireARAT_0_wen,
  output wire [4:0]    io_retireARAT_1_ard,
  output wire [5:0]    io_retireARAT_1_prd,
  output wire          io_retireARAT_1_wen,
  output wire [5:0]    io_retireFreeList_prfIdx_0,
  output wire [5:0]    io_retireFreeList_prfIdx_1,
  output wire [1:0]    io_retireFreeList_writeNum,
  output wire          io_retireFreeList_delayedFlush,
  output wire [4:0]    io_retireLSU_robIdx_0,
  output wire [4:0]    io_retireLSU_robIdx_1,
  output wire          io_retireLSU_allowRetire_0,
  output wire          io_retireLSU_allowRetire_1,
  output wire          io_wakeupMem,
  output wire          io_updateBPU_0_valid,
  output wire [31:0]   io_updateBPU_0_payload_pc,
  output wire          io_updateBPU_0_payload_isJumpInst,
  output wire          io_updateBPU_0_payload_taken,
  output wire          io_updateBPU_0_payload_predictFail,
  output wire [31:0]   io_updateBPU_0_payload_target,
  output wire          io_updateBPU_1_valid,
  output wire [31:0]   io_updateBPU_1_payload_pc,
  output wire          io_updateBPU_1_payload_isJumpInst,
  output wire          io_updateBPU_1_payload_taken,
  output wire          io_updateBPU_1_payload_predictFail,
  output wire [31:0]   io_updateBPU_1_payload_target,
  output wire          io_csrCtrl_llBitUpdate,
  output wire          io_csrCtrl_writeCSR,
  output wire          io_csrCtrl_ertn,
  output wire          io_csrCtrl_normalException,
  output wire          io_csrCtrl_tlbrException,
  output wire [31:0]   io_csrCtrl_epc,
  output wire [4:0]    io_csrCtrl_eROBIdx,
  output wire [5:0]    io_csrCtrl_eCode,
  output wire [0:0]    io_csrCtrl_eSubCode,
  input  wire [31:0]   io_csrCtrl_era,
  input  wire [31:0]   io_csrCtrl_eentry,
  input  wire [31:0]   io_csrCtrl_tlbrentry,
  output wire          io_flush,
  input  wire          io_interrupt,
  output wire [31:0]   io_redirectPC,
  output reg  [31:0]   io_commitROBEntries_0_pc,
  output reg  [4:0]    io_commitROBEntries_0_ard,
  output reg  [5:0]    io_commitROBEntries_0_prd,
  output reg  [5:0]    io_commitROBEntries_0_pprd,
  output reg  [3:0]    io_commitROBEntries_0_specialOp,
  output reg           io_commitROBEntries_0_isComplete,
  output reg  [31:0]   io_commitROBEntries_0_branchResult_targetPC,
  output reg           io_commitROBEntries_0_branchResult_branchResult,
  output reg           io_commitROBEntries_0_branchResult_predictFail,
  output reg           io_commitROBEntries_0_exceptionInfo_exception,
  output reg  [5:0]    io_commitROBEntries_0_exceptionInfo_eCode,
  output reg  [0:0]    io_commitROBEntries_0_exceptionInfo_eSubCode,
  output reg           io_commitROBEntries_0_valid,
  output reg  [31:0]   io_commitROBEntries_1_pc,
  output reg  [4:0]    io_commitROBEntries_1_ard,
  output reg  [5:0]    io_commitROBEntries_1_prd,
  output reg  [5:0]    io_commitROBEntries_1_pprd,
  output reg  [3:0]    io_commitROBEntries_1_specialOp,
  output reg           io_commitROBEntries_1_isComplete,
  output reg  [31:0]   io_commitROBEntries_1_branchResult_targetPC,
  output reg           io_commitROBEntries_1_branchResult_branchResult,
  output reg           io_commitROBEntries_1_branchResult_predictFail,
  output reg           io_commitROBEntries_1_exceptionInfo_exception,
  output reg  [5:0]    io_commitROBEntries_1_exceptionInfo_eCode,
  output reg  [0:0]    io_commitROBEntries_1_exceptionInfo_eSubCode,
  output reg           io_commitROBEntries_1_valid,
  output reg  [31:0]   io_commitROBEntries_2_pc,
  output reg  [4:0]    io_commitROBEntries_2_ard,
  output reg  [5:0]    io_commitROBEntries_2_prd,
  output reg  [5:0]    io_commitROBEntries_2_pprd,
  output reg  [3:0]    io_commitROBEntries_2_specialOp,
  output reg           io_commitROBEntries_2_isComplete,
  output reg  [31:0]   io_commitROBEntries_2_branchResult_targetPC,
  output reg           io_commitROBEntries_2_branchResult_branchResult,
  output reg           io_commitROBEntries_2_branchResult_predictFail,
  output reg           io_commitROBEntries_2_exceptionInfo_exception,
  output reg  [5:0]    io_commitROBEntries_2_exceptionInfo_eCode,
  output reg  [0:0]    io_commitROBEntries_2_exceptionInfo_eSubCode,
  output reg           io_commitROBEntries_2_valid,
  output reg  [31:0]   io_commitROBEntries_3_pc,
  output reg  [4:0]    io_commitROBEntries_3_ard,
  output reg  [5:0]    io_commitROBEntries_3_prd,
  output reg  [5:0]    io_commitROBEntries_3_pprd,
  output reg  [3:0]    io_commitROBEntries_3_specialOp,
  output reg           io_commitROBEntries_3_isComplete,
  output reg  [31:0]   io_commitROBEntries_3_branchResult_targetPC,
  output reg           io_commitROBEntries_3_branchResult_branchResult,
  output reg           io_commitROBEntries_3_branchResult_predictFail,
  output reg           io_commitROBEntries_3_exceptionInfo_exception,
  output reg  [5:0]    io_commitROBEntries_3_exceptionInfo_eCode,
  output reg  [0:0]    io_commitROBEntries_3_exceptionInfo_eSubCode,
  output reg           io_commitROBEntries_3_valid,
  output reg  [31:0]   io_commitROBEntries_4_pc,
  output reg  [4:0]    io_commitROBEntries_4_ard,
  output reg  [5:0]    io_commitROBEntries_4_prd,
  output reg  [5:0]    io_commitROBEntries_4_pprd,
  output reg  [3:0]    io_commitROBEntries_4_specialOp,
  output reg           io_commitROBEntries_4_isComplete,
  output reg  [31:0]   io_commitROBEntries_4_branchResult_targetPC,
  output reg           io_commitROBEntries_4_branchResult_branchResult,
  output reg           io_commitROBEntries_4_branchResult_predictFail,
  output reg           io_commitROBEntries_4_exceptionInfo_exception,
  output reg  [5:0]    io_commitROBEntries_4_exceptionInfo_eCode,
  output reg  [0:0]    io_commitROBEntries_4_exceptionInfo_eSubCode,
  output reg           io_commitROBEntries_4_valid,
  input  wire          aclk,
  input  wire          aresetn
);
  localparam ROBSpecialOp_nop = 4'd0;
  localparam ROBSpecialOp_bpuUpdate = 4'd1;
  localparam ROBSpecialOp_lsuAction = 4'd2;
  localparam ROBSpecialOp_ll = 4'd3;
  localparam ROBSpecialOp_writeCSR = 4'd4;
  localparam ROBSpecialOp_ertn = 4'd5;
  localparam ROBSpecialOp_idle = 4'd6;
  localparam ROBSpecialOp_readCSR = 4'd7;
  localparam ROBSpecialOp_readCNT = 4'd8;

  reg        [31:0]   _zz__zz_retirePC_0;
  reg        [5:0]    _zz__zz_noPPRDMask;
  reg        [3:0]    _zz__zz_stage_updateBPU_0_isJumpInst;
  reg                 _zz__zz_retireMask;
  reg                 _zz__zz_stage_updateBPU_0_taken;
  reg                 _zz__zz_stage_updateBPU_0_predictFail;
  reg                 _zz__zz_retireMask_1;
  reg        [5:0]    _zz__zz_normalExceptionMask;
  reg        [0:0]    _zz__zz_normalExceptionMask_1;
  reg                 _zz__zz_retireMask_2;
  reg        [1:0]    _zz_dispatchNum;
  wire       [1:0]    _zz_dispatchNum_1;
  reg        [1:0]    _zz_retireNum;
  wire       [1:0]    _zz_retireNum_1;
  reg                 _zz_stage_availROBMask;
  wire       [4:0]    _zz_stage_availROBMask_1;
  wire       [4:0]    _zz_stage_availROBMask_2;
  reg                 _zz_stage_availROBMask_3;
  wire       [4:0]    _zz_stage_availROBMask_4;
  wire       [4:0]    _zz_stage_availROBMask_5;
  reg        [31:0]   _zz__zz_retirePC_1;
  reg        [3:0]    _zz__zz_stage_updateBPU_1_isJumpInst;
  reg                 _zz__zz_retireMask_3;
  reg                 _zz__zz_stage_updateBPU_1_taken;
  reg                 _zz__zz_stage_updateBPU_1_predictFail;
  reg                 _zz__zz_retireMask_4;
  reg        [5:0]    _zz__zz_normalExceptionMask_2;
  reg        [0:0]    _zz__zz_normalExceptionMask_3;
  reg                 _zz__zz_retireMask_5;
  wire       [4:0]    _zz_tail_0;
  wire       [4:0]    _zz_tail_0_1;
  wire       [4:0]    _zz_tail_1;
  wire       [0:0]    _zz_tail_1_1;
  wire       [4:0]    _zz_tail_1_2;
  wire       [4:0]    _zz_tail_1_3;
  reg        [3:0]    _zz__zz_io_commitROBEntries_0_specialOp;
  reg        [31:0]   _zz_io_commitROBEntries_0_pc_1;
  reg        [4:0]    _zz_io_commitROBEntries_0_ard;
  reg        [5:0]    _zz_io_commitROBEntries_0_prd;
  reg        [5:0]    _zz_io_commitROBEntries_0_pprd;
  reg                 _zz_io_commitROBEntries_0_isComplete;
  reg        [31:0]   _zz_io_commitROBEntries_0_branchResult_targetPC;
  reg                 _zz_io_commitROBEntries_0_branchResult_branchResult;
  reg                 _zz_io_commitROBEntries_0_branchResult_predictFail;
  reg                 _zz_io_commitROBEntries_0_exceptionInfo_exception;
  reg        [5:0]    _zz_io_commitROBEntries_0_exceptionInfo_eCode;
  reg        [0:0]    _zz_io_commitROBEntries_0_exceptionInfo_eSubCode;
  reg                 _zz_io_commitROBEntries_0_valid;
  reg        [3:0]    _zz__zz_io_commitROBEntries_1_specialOp;
  reg        [31:0]   _zz_io_commitROBEntries_1_pc_1;
  reg        [4:0]    _zz_io_commitROBEntries_1_ard;
  reg        [5:0]    _zz_io_commitROBEntries_1_prd;
  reg        [5:0]    _zz_io_commitROBEntries_1_pprd;
  reg                 _zz_io_commitROBEntries_1_isComplete;
  reg        [31:0]   _zz_io_commitROBEntries_1_branchResult_targetPC;
  reg                 _zz_io_commitROBEntries_1_branchResult_branchResult;
  reg                 _zz_io_commitROBEntries_1_branchResult_predictFail;
  reg                 _zz_io_commitROBEntries_1_exceptionInfo_exception;
  reg        [5:0]    _zz_io_commitROBEntries_1_exceptionInfo_eCode;
  reg        [0:0]    _zz_io_commitROBEntries_1_exceptionInfo_eSubCode;
  reg                 _zz_io_commitROBEntries_1_valid;
  reg        [3:0]    _zz__zz_io_commitROBEntries_2_specialOp;
  reg        [31:0]   _zz_io_commitROBEntries_2_pc_1;
  reg        [4:0]    _zz_io_commitROBEntries_2_ard;
  reg        [5:0]    _zz_io_commitROBEntries_2_prd;
  reg        [5:0]    _zz_io_commitROBEntries_2_pprd;
  reg                 _zz_io_commitROBEntries_2_isComplete;
  reg        [31:0]   _zz_io_commitROBEntries_2_branchResult_targetPC;
  reg                 _zz_io_commitROBEntries_2_branchResult_branchResult;
  reg                 _zz_io_commitROBEntries_2_branchResult_predictFail;
  reg                 _zz_io_commitROBEntries_2_exceptionInfo_exception;
  reg        [5:0]    _zz_io_commitROBEntries_2_exceptionInfo_eCode;
  reg        [0:0]    _zz_io_commitROBEntries_2_exceptionInfo_eSubCode;
  reg                 _zz_io_commitROBEntries_2_valid;
  reg        [3:0]    _zz__zz_io_commitROBEntries_3_specialOp;
  reg        [31:0]   _zz_io_commitROBEntries_3_pc_1;
  reg        [4:0]    _zz_io_commitROBEntries_3_ard;
  reg        [5:0]    _zz_io_commitROBEntries_3_prd;
  reg        [5:0]    _zz_io_commitROBEntries_3_pprd;
  reg                 _zz_io_commitROBEntries_3_isComplete;
  reg        [31:0]   _zz_io_commitROBEntries_3_branchResult_targetPC;
  reg                 _zz_io_commitROBEntries_3_branchResult_branchResult;
  reg                 _zz_io_commitROBEntries_3_branchResult_predictFail;
  reg                 _zz_io_commitROBEntries_3_exceptionInfo_exception;
  reg        [5:0]    _zz_io_commitROBEntries_3_exceptionInfo_eCode;
  reg        [0:0]    _zz_io_commitROBEntries_3_exceptionInfo_eSubCode;
  reg                 _zz_io_commitROBEntries_3_valid;
  reg        [3:0]    _zz__zz_io_commitROBEntries_4_specialOp;
  reg        [31:0]   _zz_io_commitROBEntries_4_pc_1;
  reg        [4:0]    _zz_io_commitROBEntries_4_ard;
  reg        [5:0]    _zz_io_commitROBEntries_4_prd;
  reg        [5:0]    _zz_io_commitROBEntries_4_pprd;
  reg                 _zz_io_commitROBEntries_4_isComplete;
  reg        [31:0]   _zz_io_commitROBEntries_4_branchResult_targetPC;
  reg                 _zz_io_commitROBEntries_4_branchResult_branchResult;
  reg                 _zz_io_commitROBEntries_4_branchResult_predictFail;
  reg                 _zz_io_commitROBEntries_4_exceptionInfo_exception;
  reg        [5:0]    _zz_io_commitROBEntries_4_exceptionInfo_eCode;
  reg        [0:0]    _zz_io_commitROBEntries_4_exceptionInfo_eSubCode;
  reg                 _zz_io_commitROBEntries_4_valid;
  wire       [4:0]    _zz_head_0;
  wire       [4:0]    _zz_head_0_1;
  wire       [4:0]    _zz_head_1;
  wire       [4:0]    _zz_head_1_1;
  wire       [1:0]    _zz_noPPRDMaskMid_1_0;
  wire       [1:0]    _zz_freePRFIdxMid_1_0;
  wire       [1:0]    _zz_noPPRDMaskMid_1_1;
  wire       [1:0]    _zz_freePRFIdxMid_1_1;
  reg        [4:0]    _zz_stage_retireARAT_0_ard;
  reg        [5:0]    _zz_stage_retireARAT_0_prd;
  reg        [31:0]   _zz_retireTargetPC_0;
  reg        [4:0]    _zz_stage_retireARAT_1_ard;
  reg        [5:0]    _zz_stage_retireARAT_1_prd;
  reg        [5:0]    _zz_noPPRDMask_1;
  reg        [31:0]   _zz_retireTargetPC_1;
  reg        [1:0]    _zz_stage_freePRFNum_1;
  wire       [1:0]    _zz_stage_freePRFNum_2;
  reg        [31:0]   rob_0_pc;
  reg        [4:0]    rob_0_ard;
  reg        [5:0]    rob_0_prd;
  reg        [5:0]    rob_0_pprd;
  reg        [3:0]    rob_0_specialOp;
  reg                 rob_0_isComplete;
  reg        [31:0]   rob_0_branchResult_targetPC;
  reg                 rob_0_branchResult_branchResult;
  reg                 rob_0_branchResult_predictFail;
  reg                 rob_0_exceptionInfo_exception;
  reg        [5:0]    rob_0_exceptionInfo_eCode;
  reg        [0:0]    rob_0_exceptionInfo_eSubCode;
  reg                 rob_0_valid;
  reg        [31:0]   rob_1_pc;
  reg        [4:0]    rob_1_ard;
  reg        [5:0]    rob_1_prd;
  reg        [5:0]    rob_1_pprd;
  reg        [3:0]    rob_1_specialOp;
  reg                 rob_1_isComplete;
  reg        [31:0]   rob_1_branchResult_targetPC;
  reg                 rob_1_branchResult_branchResult;
  reg                 rob_1_branchResult_predictFail;
  reg                 rob_1_exceptionInfo_exception;
  reg        [5:0]    rob_1_exceptionInfo_eCode;
  reg        [0:0]    rob_1_exceptionInfo_eSubCode;
  reg                 rob_1_valid;
  reg        [31:0]   rob_2_pc;
  reg        [4:0]    rob_2_ard;
  reg        [5:0]    rob_2_prd;
  reg        [5:0]    rob_2_pprd;
  reg        [3:0]    rob_2_specialOp;
  reg                 rob_2_isComplete;
  reg        [31:0]   rob_2_branchResult_targetPC;
  reg                 rob_2_branchResult_branchResult;
  reg                 rob_2_branchResult_predictFail;
  reg                 rob_2_exceptionInfo_exception;
  reg        [5:0]    rob_2_exceptionInfo_eCode;
  reg        [0:0]    rob_2_exceptionInfo_eSubCode;
  reg                 rob_2_valid;
  reg        [31:0]   rob_3_pc;
  reg        [4:0]    rob_3_ard;
  reg        [5:0]    rob_3_prd;
  reg        [5:0]    rob_3_pprd;
  reg        [3:0]    rob_3_specialOp;
  reg                 rob_3_isComplete;
  reg        [31:0]   rob_3_branchResult_targetPC;
  reg                 rob_3_branchResult_branchResult;
  reg                 rob_3_branchResult_predictFail;
  reg                 rob_3_exceptionInfo_exception;
  reg        [5:0]    rob_3_exceptionInfo_eCode;
  reg        [0:0]    rob_3_exceptionInfo_eSubCode;
  reg                 rob_3_valid;
  reg        [31:0]   rob_4_pc;
  reg        [4:0]    rob_4_ard;
  reg        [5:0]    rob_4_prd;
  reg        [5:0]    rob_4_pprd;
  reg        [3:0]    rob_4_specialOp;
  reg                 rob_4_isComplete;
  reg        [31:0]   rob_4_branchResult_targetPC;
  reg                 rob_4_branchResult_branchResult;
  reg                 rob_4_branchResult_predictFail;
  reg                 rob_4_exceptionInfo_exception;
  reg        [5:0]    rob_4_exceptionInfo_eCode;
  reg        [0:0]    rob_4_exceptionInfo_eSubCode;
  reg                 rob_4_valid;
  reg        [31:0]   rob_5_pc;
  reg        [4:0]    rob_5_ard;
  reg        [5:0]    rob_5_prd;
  reg        [5:0]    rob_5_pprd;
  reg        [3:0]    rob_5_specialOp;
  reg                 rob_5_isComplete;
  reg        [31:0]   rob_5_branchResult_targetPC;
  reg                 rob_5_branchResult_branchResult;
  reg                 rob_5_branchResult_predictFail;
  reg                 rob_5_exceptionInfo_exception;
  reg        [5:0]    rob_5_exceptionInfo_eCode;
  reg        [0:0]    rob_5_exceptionInfo_eSubCode;
  reg                 rob_5_valid;
  reg        [31:0]   rob_6_pc;
  reg        [4:0]    rob_6_ard;
  reg        [5:0]    rob_6_prd;
  reg        [5:0]    rob_6_pprd;
  reg        [3:0]    rob_6_specialOp;
  reg                 rob_6_isComplete;
  reg        [31:0]   rob_6_branchResult_targetPC;
  reg                 rob_6_branchResult_branchResult;
  reg                 rob_6_branchResult_predictFail;
  reg                 rob_6_exceptionInfo_exception;
  reg        [5:0]    rob_6_exceptionInfo_eCode;
  reg        [0:0]    rob_6_exceptionInfo_eSubCode;
  reg                 rob_6_valid;
  reg        [31:0]   rob_7_pc;
  reg        [4:0]    rob_7_ard;
  reg        [5:0]    rob_7_prd;
  reg        [5:0]    rob_7_pprd;
  reg        [3:0]    rob_7_specialOp;
  reg                 rob_7_isComplete;
  reg        [31:0]   rob_7_branchResult_targetPC;
  reg                 rob_7_branchResult_branchResult;
  reg                 rob_7_branchResult_predictFail;
  reg                 rob_7_exceptionInfo_exception;
  reg        [5:0]    rob_7_exceptionInfo_eCode;
  reg        [0:0]    rob_7_exceptionInfo_eSubCode;
  reg                 rob_7_valid;
  reg        [31:0]   rob_8_pc;
  reg        [4:0]    rob_8_ard;
  reg        [5:0]    rob_8_prd;
  reg        [5:0]    rob_8_pprd;
  reg        [3:0]    rob_8_specialOp;
  reg                 rob_8_isComplete;
  reg        [31:0]   rob_8_branchResult_targetPC;
  reg                 rob_8_branchResult_branchResult;
  reg                 rob_8_branchResult_predictFail;
  reg                 rob_8_exceptionInfo_exception;
  reg        [5:0]    rob_8_exceptionInfo_eCode;
  reg        [0:0]    rob_8_exceptionInfo_eSubCode;
  reg                 rob_8_valid;
  reg        [31:0]   rob_9_pc;
  reg        [4:0]    rob_9_ard;
  reg        [5:0]    rob_9_prd;
  reg        [5:0]    rob_9_pprd;
  reg        [3:0]    rob_9_specialOp;
  reg                 rob_9_isComplete;
  reg        [31:0]   rob_9_branchResult_targetPC;
  reg                 rob_9_branchResult_branchResult;
  reg                 rob_9_branchResult_predictFail;
  reg                 rob_9_exceptionInfo_exception;
  reg        [5:0]    rob_9_exceptionInfo_eCode;
  reg        [0:0]    rob_9_exceptionInfo_eSubCode;
  reg                 rob_9_valid;
  reg        [31:0]   rob_10_pc;
  reg        [4:0]    rob_10_ard;
  reg        [5:0]    rob_10_prd;
  reg        [5:0]    rob_10_pprd;
  reg        [3:0]    rob_10_specialOp;
  reg                 rob_10_isComplete;
  reg        [31:0]   rob_10_branchResult_targetPC;
  reg                 rob_10_branchResult_branchResult;
  reg                 rob_10_branchResult_predictFail;
  reg                 rob_10_exceptionInfo_exception;
  reg        [5:0]    rob_10_exceptionInfo_eCode;
  reg        [0:0]    rob_10_exceptionInfo_eSubCode;
  reg                 rob_10_valid;
  reg        [31:0]   rob_11_pc;
  reg        [4:0]    rob_11_ard;
  reg        [5:0]    rob_11_prd;
  reg        [5:0]    rob_11_pprd;
  reg        [3:0]    rob_11_specialOp;
  reg                 rob_11_isComplete;
  reg        [31:0]   rob_11_branchResult_targetPC;
  reg                 rob_11_branchResult_branchResult;
  reg                 rob_11_branchResult_predictFail;
  reg                 rob_11_exceptionInfo_exception;
  reg        [5:0]    rob_11_exceptionInfo_eCode;
  reg        [0:0]    rob_11_exceptionInfo_eSubCode;
  reg                 rob_11_valid;
  reg        [31:0]   rob_12_pc;
  reg        [4:0]    rob_12_ard;
  reg        [5:0]    rob_12_prd;
  reg        [5:0]    rob_12_pprd;
  reg        [3:0]    rob_12_specialOp;
  reg                 rob_12_isComplete;
  reg        [31:0]   rob_12_branchResult_targetPC;
  reg                 rob_12_branchResult_branchResult;
  reg                 rob_12_branchResult_predictFail;
  reg                 rob_12_exceptionInfo_exception;
  reg        [5:0]    rob_12_exceptionInfo_eCode;
  reg        [0:0]    rob_12_exceptionInfo_eSubCode;
  reg                 rob_12_valid;
  reg        [31:0]   rob_13_pc;
  reg        [4:0]    rob_13_ard;
  reg        [5:0]    rob_13_prd;
  reg        [5:0]    rob_13_pprd;
  reg        [3:0]    rob_13_specialOp;
  reg                 rob_13_isComplete;
  reg        [31:0]   rob_13_branchResult_targetPC;
  reg                 rob_13_branchResult_branchResult;
  reg                 rob_13_branchResult_predictFail;
  reg                 rob_13_exceptionInfo_exception;
  reg        [5:0]    rob_13_exceptionInfo_eCode;
  reg        [0:0]    rob_13_exceptionInfo_eSubCode;
  reg                 rob_13_valid;
  reg        [31:0]   rob_14_pc;
  reg        [4:0]    rob_14_ard;
  reg        [5:0]    rob_14_prd;
  reg        [5:0]    rob_14_pprd;
  reg        [3:0]    rob_14_specialOp;
  reg                 rob_14_isComplete;
  reg        [31:0]   rob_14_branchResult_targetPC;
  reg                 rob_14_branchResult_branchResult;
  reg                 rob_14_branchResult_predictFail;
  reg                 rob_14_exceptionInfo_exception;
  reg        [5:0]    rob_14_exceptionInfo_eCode;
  reg        [0:0]    rob_14_exceptionInfo_eSubCode;
  reg                 rob_14_valid;
  reg        [31:0]   rob_15_pc;
  reg        [4:0]    rob_15_ard;
  reg        [5:0]    rob_15_prd;
  reg        [5:0]    rob_15_pprd;
  reg        [3:0]    rob_15_specialOp;
  reg                 rob_15_isComplete;
  reg        [31:0]   rob_15_branchResult_targetPC;
  reg                 rob_15_branchResult_branchResult;
  reg                 rob_15_branchResult_predictFail;
  reg                 rob_15_exceptionInfo_exception;
  reg        [5:0]    rob_15_exceptionInfo_eCode;
  reg        [0:0]    rob_15_exceptionInfo_eSubCode;
  reg                 rob_15_valid;
  reg        [31:0]   rob_16_pc;
  reg        [4:0]    rob_16_ard;
  reg        [5:0]    rob_16_prd;
  reg        [5:0]    rob_16_pprd;
  reg        [3:0]    rob_16_specialOp;
  reg                 rob_16_isComplete;
  reg        [31:0]   rob_16_branchResult_targetPC;
  reg                 rob_16_branchResult_branchResult;
  reg                 rob_16_branchResult_predictFail;
  reg                 rob_16_exceptionInfo_exception;
  reg        [5:0]    rob_16_exceptionInfo_eCode;
  reg        [0:0]    rob_16_exceptionInfo_eSubCode;
  reg                 rob_16_valid;
  reg        [31:0]   rob_17_pc;
  reg        [4:0]    rob_17_ard;
  reg        [5:0]    rob_17_prd;
  reg        [5:0]    rob_17_pprd;
  reg        [3:0]    rob_17_specialOp;
  reg                 rob_17_isComplete;
  reg        [31:0]   rob_17_branchResult_targetPC;
  reg                 rob_17_branchResult_branchResult;
  reg                 rob_17_branchResult_predictFail;
  reg                 rob_17_exceptionInfo_exception;
  reg        [5:0]    rob_17_exceptionInfo_eCode;
  reg        [0:0]    rob_17_exceptionInfo_eSubCode;
  reg                 rob_17_valid;
  reg        [31:0]   rob_18_pc;
  reg        [4:0]    rob_18_ard;
  reg        [5:0]    rob_18_prd;
  reg        [5:0]    rob_18_pprd;
  reg        [3:0]    rob_18_specialOp;
  reg                 rob_18_isComplete;
  reg        [31:0]   rob_18_branchResult_targetPC;
  reg                 rob_18_branchResult_branchResult;
  reg                 rob_18_branchResult_predictFail;
  reg                 rob_18_exceptionInfo_exception;
  reg        [5:0]    rob_18_exceptionInfo_eCode;
  reg        [0:0]    rob_18_exceptionInfo_eSubCode;
  reg                 rob_18_valid;
  reg        [31:0]   rob_19_pc;
  reg        [4:0]    rob_19_ard;
  reg        [5:0]    rob_19_prd;
  reg        [5:0]    rob_19_pprd;
  reg        [3:0]    rob_19_specialOp;
  reg                 rob_19_isComplete;
  reg        [31:0]   rob_19_branchResult_targetPC;
  reg                 rob_19_branchResult_branchResult;
  reg                 rob_19_branchResult_predictFail;
  reg                 rob_19_exceptionInfo_exception;
  reg        [5:0]    rob_19_exceptionInfo_eCode;
  reg        [0:0]    rob_19_exceptionInfo_eSubCode;
  reg                 rob_19_valid;
  reg        [31:0]   rob_20_pc;
  reg        [4:0]    rob_20_ard;
  reg        [5:0]    rob_20_prd;
  reg        [5:0]    rob_20_pprd;
  reg        [3:0]    rob_20_specialOp;
  reg                 rob_20_isComplete;
  reg        [31:0]   rob_20_branchResult_targetPC;
  reg                 rob_20_branchResult_branchResult;
  reg                 rob_20_branchResult_predictFail;
  reg                 rob_20_exceptionInfo_exception;
  reg        [5:0]    rob_20_exceptionInfo_eCode;
  reg        [0:0]    rob_20_exceptionInfo_eSubCode;
  reg                 rob_20_valid;
  reg        [31:0]   rob_21_pc;
  reg        [4:0]    rob_21_ard;
  reg        [5:0]    rob_21_prd;
  reg        [5:0]    rob_21_pprd;
  reg        [3:0]    rob_21_specialOp;
  reg                 rob_21_isComplete;
  reg        [31:0]   rob_21_branchResult_targetPC;
  reg                 rob_21_branchResult_branchResult;
  reg                 rob_21_branchResult_predictFail;
  reg                 rob_21_exceptionInfo_exception;
  reg        [5:0]    rob_21_exceptionInfo_eCode;
  reg        [0:0]    rob_21_exceptionInfo_eSubCode;
  reg                 rob_21_valid;
  reg        [31:0]   rob_22_pc;
  reg        [4:0]    rob_22_ard;
  reg        [5:0]    rob_22_prd;
  reg        [5:0]    rob_22_pprd;
  reg        [3:0]    rob_22_specialOp;
  reg                 rob_22_isComplete;
  reg        [31:0]   rob_22_branchResult_targetPC;
  reg                 rob_22_branchResult_branchResult;
  reg                 rob_22_branchResult_predictFail;
  reg                 rob_22_exceptionInfo_exception;
  reg        [5:0]    rob_22_exceptionInfo_eCode;
  reg        [0:0]    rob_22_exceptionInfo_eSubCode;
  reg                 rob_22_valid;
  reg        [31:0]   rob_23_pc;
  reg        [4:0]    rob_23_ard;
  reg        [5:0]    rob_23_prd;
  reg        [5:0]    rob_23_pprd;
  reg        [3:0]    rob_23_specialOp;
  reg                 rob_23_isComplete;
  reg        [31:0]   rob_23_branchResult_targetPC;
  reg                 rob_23_branchResult_branchResult;
  reg                 rob_23_branchResult_predictFail;
  reg                 rob_23_exceptionInfo_exception;
  reg        [5:0]    rob_23_exceptionInfo_eCode;
  reg        [0:0]    rob_23_exceptionInfo_eSubCode;
  reg                 rob_23_valid;
  reg        [31:0]   rob_24_pc;
  reg        [4:0]    rob_24_ard;
  reg        [5:0]    rob_24_prd;
  reg        [5:0]    rob_24_pprd;
  reg        [3:0]    rob_24_specialOp;
  reg                 rob_24_isComplete;
  reg        [31:0]   rob_24_branchResult_targetPC;
  reg                 rob_24_branchResult_branchResult;
  reg                 rob_24_branchResult_predictFail;
  reg                 rob_24_exceptionInfo_exception;
  reg        [5:0]    rob_24_exceptionInfo_eCode;
  reg        [0:0]    rob_24_exceptionInfo_eSubCode;
  reg                 rob_24_valid;
  reg        [31:0]   rob_25_pc;
  reg        [4:0]    rob_25_ard;
  reg        [5:0]    rob_25_prd;
  reg        [5:0]    rob_25_pprd;
  reg        [3:0]    rob_25_specialOp;
  reg                 rob_25_isComplete;
  reg        [31:0]   rob_25_branchResult_targetPC;
  reg                 rob_25_branchResult_branchResult;
  reg                 rob_25_branchResult_predictFail;
  reg                 rob_25_exceptionInfo_exception;
  reg        [5:0]    rob_25_exceptionInfo_eCode;
  reg        [0:0]    rob_25_exceptionInfo_eSubCode;
  reg                 rob_25_valid;
  reg        [31:0]   rob_26_pc;
  reg        [4:0]    rob_26_ard;
  reg        [5:0]    rob_26_prd;
  reg        [5:0]    rob_26_pprd;
  reg        [3:0]    rob_26_specialOp;
  reg                 rob_26_isComplete;
  reg        [31:0]   rob_26_branchResult_targetPC;
  reg                 rob_26_branchResult_branchResult;
  reg                 rob_26_branchResult_predictFail;
  reg                 rob_26_exceptionInfo_exception;
  reg        [5:0]    rob_26_exceptionInfo_eCode;
  reg        [0:0]    rob_26_exceptionInfo_eSubCode;
  reg                 rob_26_valid;
  reg        [31:0]   rob_27_pc;
  reg        [4:0]    rob_27_ard;
  reg        [5:0]    rob_27_prd;
  reg        [5:0]    rob_27_pprd;
  reg        [3:0]    rob_27_specialOp;
  reg                 rob_27_isComplete;
  reg        [31:0]   rob_27_branchResult_targetPC;
  reg                 rob_27_branchResult_branchResult;
  reg                 rob_27_branchResult_predictFail;
  reg                 rob_27_exceptionInfo_exception;
  reg        [5:0]    rob_27_exceptionInfo_eCode;
  reg        [0:0]    rob_27_exceptionInfo_eSubCode;
  reg                 rob_27_valid;
  reg        [31:0]   rob_28_pc;
  reg        [4:0]    rob_28_ard;
  reg        [5:0]    rob_28_prd;
  reg        [5:0]    rob_28_pprd;
  reg        [3:0]    rob_28_specialOp;
  reg                 rob_28_isComplete;
  reg        [31:0]   rob_28_branchResult_targetPC;
  reg                 rob_28_branchResult_branchResult;
  reg                 rob_28_branchResult_predictFail;
  reg                 rob_28_exceptionInfo_exception;
  reg        [5:0]    rob_28_exceptionInfo_eCode;
  reg        [0:0]    rob_28_exceptionInfo_eSubCode;
  reg                 rob_28_valid;
  reg        [31:0]   rob_29_pc;
  reg        [4:0]    rob_29_ard;
  reg        [5:0]    rob_29_prd;
  reg        [5:0]    rob_29_pprd;
  reg        [3:0]    rob_29_specialOp;
  reg                 rob_29_isComplete;
  reg        [31:0]   rob_29_branchResult_targetPC;
  reg                 rob_29_branchResult_branchResult;
  reg                 rob_29_branchResult_predictFail;
  reg                 rob_29_exceptionInfo_exception;
  reg        [5:0]    rob_29_exceptionInfo_eCode;
  reg        [0:0]    rob_29_exceptionInfo_eSubCode;
  reg                 rob_29_valid;
  reg        [31:0]   rob_30_pc;
  reg        [4:0]    rob_30_ard;
  reg        [5:0]    rob_30_prd;
  reg        [5:0]    rob_30_pprd;
  reg        [3:0]    rob_30_specialOp;
  reg                 rob_30_isComplete;
  reg        [31:0]   rob_30_branchResult_targetPC;
  reg                 rob_30_branchResult_branchResult;
  reg                 rob_30_branchResult_predictFail;
  reg                 rob_30_exceptionInfo_exception;
  reg        [5:0]    rob_30_exceptionInfo_eCode;
  reg        [0:0]    rob_30_exceptionInfo_eSubCode;
  reg                 rob_30_valid;
  reg        [31:0]   rob_31_pc;
  reg        [4:0]    rob_31_ard;
  reg        [5:0]    rob_31_prd;
  reg        [5:0]    rob_31_pprd;
  reg        [3:0]    rob_31_specialOp;
  reg                 rob_31_isComplete;
  reg        [31:0]   rob_31_branchResult_targetPC;
  reg                 rob_31_branchResult_branchResult;
  reg                 rob_31_branchResult_predictFail;
  reg                 rob_31_exceptionInfo_exception;
  reg        [5:0]    rob_31_exceptionInfo_eCode;
  reg        [0:0]    rob_31_exceptionInfo_eSubCode;
  reg                 rob_31_valid;
  reg        [4:0]    head_0;
  reg        [4:0]    head_1;
  reg        [4:0]    tail_0;
  reg        [4:0]    tail_1;
  reg        [1:0]    stage_availROBMask;
  wire       [4:0]    stage_retireARAT_0_ard;
  wire       [5:0]    stage_retireARAT_0_prd;
  wire                stage_retireARAT_0_wen;
  wire       [4:0]    stage_retireARAT_1_ard;
  wire       [5:0]    stage_retireARAT_1_prd;
  wire                stage_retireARAT_1_wen;
  wire       [5:0]    stage_freePRFIdx_0;
  wire       [5:0]    stage_freePRFIdx_1;
  wire       [1:0]    stage_freePRFNum;
  wire       [4:0]    stage_retireROBIdx_0;
  wire       [4:0]    stage_retireROBIdx_1;
  wire                stage_retireEn_0;
  wire                stage_retireEn_1;
  wire                stage_wakeupMem;
  wire                stage_retireLLBitUpdate;
  wire                stage_retireWriteCSR;
  wire                stage_retireERTN;
  wire                stage_retireNormalException;
  wire                stage_retireTLBRException;
  wire       [31:0]   stage_retireEPC;
  wire       [4:0]    stage_retireEROBIdx;
  wire       [5:0]    stage_retireECode;
  wire       [0:0]    stage_retireESubCode;
  wire       [31:0]   stage_updateBPU_0_pc;
  wire                stage_updateBPU_0_isJumpInst;
  wire                stage_updateBPU_0_taken;
  wire                stage_updateBPU_0_predictFail;
  wire       [31:0]   stage_updateBPU_0_target;
  wire       [31:0]   stage_updateBPU_1_pc;
  wire                stage_updateBPU_1_isJumpInst;
  wire                stage_updateBPU_1_taken;
  wire                stage_updateBPU_1_predictFail;
  wire       [31:0]   stage_updateBPU_1_target;
  wire                stage_flush;
  wire       [31:0]   stage_redirectPC;
  reg        [1:0]    retireMask;
  reg        [1:0]    inhibitNextRetireMask;
  reg        [1:0]    flushMask;
  wire                flush;
  wire       [31:0]   _zz_retirePC_0;
  wire       [5:0]    _zz_noPPRDMask;
  wire       [3:0]    _zz_stage_updateBPU_0_isJumpInst;
  wire                _zz_retireMask;
  wire                _zz_stage_updateBPU_0_taken;
  wire                _zz_stage_updateBPU_0_predictFail;
  wire                _zz_retireMask_1;
  wire       [5:0]    _zz_normalExceptionMask;
  wire       [0:0]    _zz_normalExceptionMask_1;
  wire                _zz_retireMask_2;
  wire                idleEn;
  wire       [1:0]    dispatchNum;
  wire       [1:0]    retireNum;
  wire       [31:0]   _zz_retirePC_1;
  wire       [3:0]    _zz_stage_updateBPU_1_isJumpInst;
  wire                _zz_retireMask_3;
  wire                _zz_stage_updateBPU_1_taken;
  wire                _zz_stage_updateBPU_1_predictFail;
  wire                _zz_retireMask_4;
  wire       [5:0]    _zz_normalExceptionMask_2;
  wire       [0:0]    _zz_normalExceptionMask_3;
  wire                _zz_retireMask_5;
  reg        [1:0]    _zz_rob_0_valid;
  reg        [4:0]    _zz_rob_0_isComplete;
  reg        [1:0]    _zz_rob_0_isComplete_1;
  reg        [1:0]    _zz_rob_1_valid;
  reg        [4:0]    _zz_rob_1_isComplete;
  reg        [1:0]    _zz_rob_1_isComplete_1;
  reg        [1:0]    _zz_rob_2_valid;
  reg        [4:0]    _zz_rob_2_isComplete;
  reg        [1:0]    _zz_rob_2_isComplete_1;
  reg        [1:0]    _zz_rob_3_valid;
  reg        [4:0]    _zz_rob_3_isComplete;
  reg        [1:0]    _zz_rob_3_isComplete_1;
  reg        [1:0]    _zz_rob_4_valid;
  reg        [4:0]    _zz_rob_4_isComplete;
  reg        [1:0]    _zz_rob_4_isComplete_1;
  reg        [1:0]    _zz_rob_5_valid;
  reg        [4:0]    _zz_rob_5_isComplete;
  reg        [1:0]    _zz_rob_5_isComplete_1;
  reg        [1:0]    _zz_rob_6_valid;
  reg        [4:0]    _zz_rob_6_isComplete;
  reg        [1:0]    _zz_rob_6_isComplete_1;
  reg        [1:0]    _zz_rob_7_valid;
  reg        [4:0]    _zz_rob_7_isComplete;
  reg        [1:0]    _zz_rob_7_isComplete_1;
  reg        [1:0]    _zz_rob_8_valid;
  reg        [4:0]    _zz_rob_8_isComplete;
  reg        [1:0]    _zz_rob_8_isComplete_1;
  reg        [1:0]    _zz_rob_9_valid;
  reg        [4:0]    _zz_rob_9_isComplete;
  reg        [1:0]    _zz_rob_9_isComplete_1;
  reg        [1:0]    _zz_rob_10_valid;
  reg        [4:0]    _zz_rob_10_isComplete;
  reg        [1:0]    _zz_rob_10_isComplete_1;
  reg        [1:0]    _zz_rob_11_valid;
  reg        [4:0]    _zz_rob_11_isComplete;
  reg        [1:0]    _zz_rob_11_isComplete_1;
  reg        [1:0]    _zz_rob_12_valid;
  reg        [4:0]    _zz_rob_12_isComplete;
  reg        [1:0]    _zz_rob_12_isComplete_1;
  reg        [1:0]    _zz_rob_13_valid;
  reg        [4:0]    _zz_rob_13_isComplete;
  reg        [1:0]    _zz_rob_13_isComplete_1;
  reg        [1:0]    _zz_rob_14_valid;
  reg        [4:0]    _zz_rob_14_isComplete;
  reg        [1:0]    _zz_rob_14_isComplete_1;
  reg        [1:0]    _zz_rob_15_valid;
  reg        [4:0]    _zz_rob_15_isComplete;
  reg        [1:0]    _zz_rob_15_isComplete_1;
  reg        [1:0]    _zz_rob_16_valid;
  reg        [4:0]    _zz_rob_16_isComplete;
  reg        [1:0]    _zz_rob_16_isComplete_1;
  reg        [1:0]    _zz_rob_17_valid;
  reg        [4:0]    _zz_rob_17_isComplete;
  reg        [1:0]    _zz_rob_17_isComplete_1;
  reg        [1:0]    _zz_rob_18_valid;
  reg        [4:0]    _zz_rob_18_isComplete;
  reg        [1:0]    _zz_rob_18_isComplete_1;
  reg        [1:0]    _zz_rob_19_valid;
  reg        [4:0]    _zz_rob_19_isComplete;
  reg        [1:0]    _zz_rob_19_isComplete_1;
  reg        [1:0]    _zz_rob_20_valid;
  reg        [4:0]    _zz_rob_20_isComplete;
  reg        [1:0]    _zz_rob_20_isComplete_1;
  reg        [1:0]    _zz_rob_21_valid;
  reg        [4:0]    _zz_rob_21_isComplete;
  reg        [1:0]    _zz_rob_21_isComplete_1;
  reg        [1:0]    _zz_rob_22_valid;
  reg        [4:0]    _zz_rob_22_isComplete;
  reg        [1:0]    _zz_rob_22_isComplete_1;
  reg        [1:0]    _zz_rob_23_valid;
  reg        [4:0]    _zz_rob_23_isComplete;
  reg        [1:0]    _zz_rob_23_isComplete_1;
  reg        [1:0]    _zz_rob_24_valid;
  reg        [4:0]    _zz_rob_24_isComplete;
  reg        [1:0]    _zz_rob_24_isComplete_1;
  reg        [1:0]    _zz_rob_25_valid;
  reg        [4:0]    _zz_rob_25_isComplete;
  reg        [1:0]    _zz_rob_25_isComplete_1;
  reg        [1:0]    _zz_rob_26_valid;
  reg        [4:0]    _zz_rob_26_isComplete;
  reg        [1:0]    _zz_rob_26_isComplete_1;
  reg        [1:0]    _zz_rob_27_valid;
  reg        [4:0]    _zz_rob_27_isComplete;
  reg        [1:0]    _zz_rob_27_isComplete_1;
  reg        [1:0]    _zz_rob_28_valid;
  reg        [4:0]    _zz_rob_28_isComplete;
  reg        [1:0]    _zz_rob_28_isComplete_1;
  reg        [1:0]    _zz_rob_29_valid;
  reg        [4:0]    _zz_rob_29_isComplete;
  reg        [1:0]    _zz_rob_29_isComplete_1;
  reg        [1:0]    _zz_rob_30_valid;
  reg        [4:0]    _zz_rob_30_isComplete;
  reg        [1:0]    _zz_rob_30_isComplete_1;
  reg        [1:0]    _zz_rob_31_valid;
  reg        [4:0]    _zz_rob_31_isComplete;
  reg        [1:0]    _zz_rob_31_isComplete_1;
  wire                when_ROB_l76;
  wire       [31:0]   _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                when_ROB_l76_1;
  wire       [31:0]   _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire       [31:0]   _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire                _zz_70;
  wire                _zz_71;
  wire                _zz_72;
  wire                _zz_73;
  wire                _zz_74;
  wire                _zz_75;
  wire                _zz_76;
  wire                _zz_77;
  wire                _zz_78;
  wire                _zz_79;
  wire                _zz_80;
  wire                _zz_81;
  wire                _zz_82;
  wire                _zz_83;
  wire                _zz_84;
  wire                _zz_85;
  wire                _zz_86;
  wire                _zz_87;
  wire                _zz_88;
  wire                _zz_89;
  wire                _zz_90;
  wire                _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire                _zz_94;
  wire                _zz_95;
  wire                _zz_96;
  wire                _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire       [31:0]   _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire                _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire                _zz_106;
  wire                _zz_107;
  wire                _zz_108;
  wire                _zz_109;
  wire                _zz_110;
  wire                _zz_111;
  wire                _zz_112;
  wire                _zz_113;
  wire                _zz_114;
  wire                _zz_115;
  wire                _zz_116;
  wire                _zz_117;
  wire                _zz_118;
  wire                _zz_119;
  wire                _zz_120;
  wire                _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire                _zz_124;
  wire                _zz_125;
  wire                _zz_126;
  wire                _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire                _zz_130;
  wire                _zz_131;
  wire                _zz_132;
  wire       [4:0]    _zz_io_commitROBEntries_0_pc;
  wire       [3:0]    _zz_io_commitROBEntries_0_specialOp;
  wire       [31:0]   _zz_133;
  wire                _zz_134;
  wire                _zz_135;
  wire                _zz_136;
  wire                _zz_137;
  wire                _zz_138;
  wire                _zz_139;
  wire                _zz_140;
  wire                _zz_141;
  wire                _zz_142;
  wire                _zz_143;
  wire                _zz_144;
  wire                _zz_145;
  wire                _zz_146;
  wire                _zz_147;
  wire                _zz_148;
  wire                _zz_149;
  wire                _zz_150;
  wire                _zz_151;
  wire                _zz_152;
  wire                _zz_153;
  wire                _zz_154;
  wire                _zz_155;
  wire                _zz_156;
  wire                _zz_157;
  wire                _zz_158;
  wire                _zz_159;
  wire                _zz_160;
  wire                _zz_161;
  wire                _zz_162;
  wire                _zz_163;
  wire                _zz_164;
  wire                _zz_165;
  wire       [31:0]   _zz_166;
  wire                _zz_167;
  wire                _zz_168;
  wire                _zz_169;
  wire                _zz_170;
  wire                _zz_171;
  wire                _zz_172;
  wire                _zz_173;
  wire                _zz_174;
  wire                _zz_175;
  wire                _zz_176;
  wire                _zz_177;
  wire                _zz_178;
  wire                _zz_179;
  wire                _zz_180;
  wire                _zz_181;
  wire                _zz_182;
  wire                _zz_183;
  wire                _zz_184;
  wire                _zz_185;
  wire                _zz_186;
  wire                _zz_187;
  wire                _zz_188;
  wire                _zz_189;
  wire                _zz_190;
  wire                _zz_191;
  wire                _zz_192;
  wire                _zz_193;
  wire                _zz_194;
  wire                _zz_195;
  wire                _zz_196;
  wire                _zz_197;
  wire                _zz_198;
  wire       [4:0]    _zz_io_commitROBEntries_1_pc;
  wire       [3:0]    _zz_io_commitROBEntries_1_specialOp;
  wire       [31:0]   _zz_199;
  wire                _zz_200;
  wire                _zz_201;
  wire                _zz_202;
  wire                _zz_203;
  wire                _zz_204;
  wire                _zz_205;
  wire                _zz_206;
  wire                _zz_207;
  wire                _zz_208;
  wire                _zz_209;
  wire                _zz_210;
  wire                _zz_211;
  wire                _zz_212;
  wire                _zz_213;
  wire                _zz_214;
  wire                _zz_215;
  wire                _zz_216;
  wire                _zz_217;
  wire                _zz_218;
  wire                _zz_219;
  wire                _zz_220;
  wire                _zz_221;
  wire                _zz_222;
  wire                _zz_223;
  wire                _zz_224;
  wire                _zz_225;
  wire                _zz_226;
  wire                _zz_227;
  wire                _zz_228;
  wire                _zz_229;
  wire                _zz_230;
  wire                _zz_231;
  wire       [31:0]   _zz_232;
  wire                _zz_233;
  wire                _zz_234;
  wire                _zz_235;
  wire                _zz_236;
  wire                _zz_237;
  wire                _zz_238;
  wire                _zz_239;
  wire                _zz_240;
  wire                _zz_241;
  wire                _zz_242;
  wire                _zz_243;
  wire                _zz_244;
  wire                _zz_245;
  wire                _zz_246;
  wire                _zz_247;
  wire                _zz_248;
  wire                _zz_249;
  wire                _zz_250;
  wire                _zz_251;
  wire                _zz_252;
  wire                _zz_253;
  wire                _zz_254;
  wire                _zz_255;
  wire                _zz_256;
  wire                _zz_257;
  wire                _zz_258;
  wire                _zz_259;
  wire                _zz_260;
  wire                _zz_261;
  wire                _zz_262;
  wire                _zz_263;
  wire                _zz_264;
  wire       [4:0]    _zz_io_commitROBEntries_2_pc;
  wire       [3:0]    _zz_io_commitROBEntries_2_specialOp;
  wire       [31:0]   _zz_265;
  wire                _zz_266;
  wire                _zz_267;
  wire                _zz_268;
  wire                _zz_269;
  wire                _zz_270;
  wire                _zz_271;
  wire                _zz_272;
  wire                _zz_273;
  wire                _zz_274;
  wire                _zz_275;
  wire                _zz_276;
  wire                _zz_277;
  wire                _zz_278;
  wire                _zz_279;
  wire                _zz_280;
  wire                _zz_281;
  wire                _zz_282;
  wire                _zz_283;
  wire                _zz_284;
  wire                _zz_285;
  wire                _zz_286;
  wire                _zz_287;
  wire                _zz_288;
  wire                _zz_289;
  wire                _zz_290;
  wire                _zz_291;
  wire                _zz_292;
  wire                _zz_293;
  wire                _zz_294;
  wire                _zz_295;
  wire                _zz_296;
  wire                _zz_297;
  wire       [31:0]   _zz_298;
  wire                _zz_299;
  wire                _zz_300;
  wire                _zz_301;
  wire                _zz_302;
  wire                _zz_303;
  wire                _zz_304;
  wire                _zz_305;
  wire                _zz_306;
  wire                _zz_307;
  wire                _zz_308;
  wire                _zz_309;
  wire                _zz_310;
  wire                _zz_311;
  wire                _zz_312;
  wire                _zz_313;
  wire                _zz_314;
  wire                _zz_315;
  wire                _zz_316;
  wire                _zz_317;
  wire                _zz_318;
  wire                _zz_319;
  wire                _zz_320;
  wire                _zz_321;
  wire                _zz_322;
  wire                _zz_323;
  wire                _zz_324;
  wire                _zz_325;
  wire                _zz_326;
  wire                _zz_327;
  wire                _zz_328;
  wire                _zz_329;
  wire                _zz_330;
  wire       [4:0]    _zz_io_commitROBEntries_3_pc;
  wire       [3:0]    _zz_io_commitROBEntries_3_specialOp;
  wire       [31:0]   _zz_331;
  wire                _zz_332;
  wire                _zz_333;
  wire                _zz_334;
  wire                _zz_335;
  wire                _zz_336;
  wire                _zz_337;
  wire                _zz_338;
  wire                _zz_339;
  wire                _zz_340;
  wire                _zz_341;
  wire                _zz_342;
  wire                _zz_343;
  wire                _zz_344;
  wire                _zz_345;
  wire                _zz_346;
  wire                _zz_347;
  wire                _zz_348;
  wire                _zz_349;
  wire                _zz_350;
  wire                _zz_351;
  wire                _zz_352;
  wire                _zz_353;
  wire                _zz_354;
  wire                _zz_355;
  wire                _zz_356;
  wire                _zz_357;
  wire                _zz_358;
  wire                _zz_359;
  wire                _zz_360;
  wire                _zz_361;
  wire                _zz_362;
  wire                _zz_363;
  wire       [31:0]   _zz_364;
  wire                _zz_365;
  wire                _zz_366;
  wire                _zz_367;
  wire                _zz_368;
  wire                _zz_369;
  wire                _zz_370;
  wire                _zz_371;
  wire                _zz_372;
  wire                _zz_373;
  wire                _zz_374;
  wire                _zz_375;
  wire                _zz_376;
  wire                _zz_377;
  wire                _zz_378;
  wire                _zz_379;
  wire                _zz_380;
  wire                _zz_381;
  wire                _zz_382;
  wire                _zz_383;
  wire                _zz_384;
  wire                _zz_385;
  wire                _zz_386;
  wire                _zz_387;
  wire                _zz_388;
  wire                _zz_389;
  wire                _zz_390;
  wire                _zz_391;
  wire                _zz_392;
  wire                _zz_393;
  wire                _zz_394;
  wire                _zz_395;
  wire                _zz_396;
  wire       [4:0]    _zz_io_commitROBEntries_4_pc;
  wire       [3:0]    _zz_io_commitROBEntries_4_specialOp;
  reg                 delayedFlush;
  reg        [1:0]    noPPRDMask;
  reg        [1:0]    lsuActionMask;
  reg        [1:0]    llMask;
  reg        [1:0]    writeCSRMask;
  reg        [1:0]    ertnMask;
  reg        [1:0]    normalExceptionMask;
  reg        [1:0]    tlbrExceptionMask;
  reg        [1:0]    falseTakenMask;
  wire       [31:0]   retirePC_0;
  wire       [31:0]   retirePC_1;
  wire       [4:0]    retireEROBIdx_0;
  wire       [4:0]    retireEROBIdx_1;
  wire       [5:0]    retireECode_0;
  wire       [5:0]    retireECode_1;
  wire       [0:0]    retireESubCode_0;
  wire       [0:0]    retireESubCode_1;
  wire       [31:0]   retireSNPC_0;
  wire       [31:0]   retireSNPC_1;
  wire       [31:0]   retireTargetPC_0;
  wire       [31:0]   retireTargetPC_1;
  wire                _zz_retireEPC;
  wire       [31:0]   retireEPC;
  wire       [4:0]    retireRealEROBIdx;
  wire       [5:0]    retireRealECode;
  wire       [0:0]    retireRealESubCode;
  wire                ertn;
  wire                normalException;
  wire                tlbrException;
  wire                falseTaken;
  wire       [31:0]   snpc;
  wire       [31:0]   targetPC;
  wire                noPPRDMaskMid_0_0;
  wire                noPPRDMaskMid_0_1;
  wire                noPPRDMaskMid_1_0;
  wire                noPPRDMaskMid_1_1;
  wire       [5:0]    freePRFIdxMid_0_0;
  wire       [5:0]    freePRFIdxMid_0_1;
  wire       [5:0]    freePRFIdxMid_1_0;
  wire       [5:0]    freePRFIdxMid_1_1;
  wire       [1:0]    _zz_stage_freePRFNum;
  reg        [1:0]    stageReg_availROBMask;
  reg        [4:0]    stageReg_retireARAT_0_ard;
  reg        [5:0]    stageReg_retireARAT_0_prd;
  reg                 stageReg_retireARAT_0_wen;
  reg        [4:0]    stageReg_retireARAT_1_ard;
  reg        [5:0]    stageReg_retireARAT_1_prd;
  reg                 stageReg_retireARAT_1_wen;
  reg        [5:0]    stageReg_freePRFIdx_0;
  reg        [5:0]    stageReg_freePRFIdx_1;
  reg        [1:0]    stageReg_freePRFNum;
  reg        [4:0]    stageReg_retireROBIdx_0;
  reg        [4:0]    stageReg_retireROBIdx_1;
  reg                 stageReg_retireEn_0;
  reg                 stageReg_retireEn_1;
  reg                 stageReg_wakeupMem;
  reg                 stageReg_retireLLBitUpdate;
  reg                 stageReg_retireWriteCSR;
  reg                 stageReg_retireERTN;
  reg                 stageReg_retireNormalException;
  reg                 stageReg_retireTLBRException;
  reg        [31:0]   stageReg_retireEPC;
  reg        [4:0]    stageReg_retireEROBIdx;
  reg        [5:0]    stageReg_retireECode;
  reg        [0:0]    stageReg_retireESubCode;
  reg        [31:0]   stageReg_updateBPU_0_pc;
  reg                 stageReg_updateBPU_0_isJumpInst;
  reg                 stageReg_updateBPU_0_taken;
  reg                 stageReg_updateBPU_0_predictFail;
  reg        [31:0]   stageReg_updateBPU_0_target;
  reg        [31:0]   stageReg_updateBPU_1_pc;
  reg                 stageReg_updateBPU_1_isJumpInst;
  reg                 stageReg_updateBPU_1_taken;
  reg                 stageReg_updateBPU_1_predictFail;
  reg        [31:0]   stageReg_updateBPU_1_target;
  reg                 stageReg_flush;
  reg        [31:0]   stageReg_redirectPC;
  `ifndef SYNTHESIS
  reg [71:0] io_dispatch_specialOp_0_string;
  reg [71:0] io_dispatch_specialOp_1_string;
  reg [71:0] io_commitROBEntries_0_specialOp_string;
  reg [71:0] io_commitROBEntries_1_specialOp_string;
  reg [71:0] io_commitROBEntries_2_specialOp_string;
  reg [71:0] io_commitROBEntries_3_specialOp_string;
  reg [71:0] io_commitROBEntries_4_specialOp_string;
  reg [71:0] rob_0_specialOp_string;
  reg [71:0] rob_1_specialOp_string;
  reg [71:0] rob_2_specialOp_string;
  reg [71:0] rob_3_specialOp_string;
  reg [71:0] rob_4_specialOp_string;
  reg [71:0] rob_5_specialOp_string;
  reg [71:0] rob_6_specialOp_string;
  reg [71:0] rob_7_specialOp_string;
  reg [71:0] rob_8_specialOp_string;
  reg [71:0] rob_9_specialOp_string;
  reg [71:0] rob_10_specialOp_string;
  reg [71:0] rob_11_specialOp_string;
  reg [71:0] rob_12_specialOp_string;
  reg [71:0] rob_13_specialOp_string;
  reg [71:0] rob_14_specialOp_string;
  reg [71:0] rob_15_specialOp_string;
  reg [71:0] rob_16_specialOp_string;
  reg [71:0] rob_17_specialOp_string;
  reg [71:0] rob_18_specialOp_string;
  reg [71:0] rob_19_specialOp_string;
  reg [71:0] rob_20_specialOp_string;
  reg [71:0] rob_21_specialOp_string;
  reg [71:0] rob_22_specialOp_string;
  reg [71:0] rob_23_specialOp_string;
  reg [71:0] rob_24_specialOp_string;
  reg [71:0] rob_25_specialOp_string;
  reg [71:0] rob_26_specialOp_string;
  reg [71:0] rob_27_specialOp_string;
  reg [71:0] rob_28_specialOp_string;
  reg [71:0] rob_29_specialOp_string;
  reg [71:0] rob_30_specialOp_string;
  reg [71:0] rob_31_specialOp_string;
  reg [71:0] _zz_stage_updateBPU_0_isJumpInst_string;
  reg [71:0] _zz_stage_updateBPU_1_isJumpInst_string;
  reg [71:0] _zz_io_commitROBEntries_0_specialOp_string;
  reg [71:0] _zz_io_commitROBEntries_1_specialOp_string;
  reg [71:0] _zz_io_commitROBEntries_2_specialOp_string;
  reg [71:0] _zz_io_commitROBEntries_3_specialOp_string;
  reg [71:0] _zz_io_commitROBEntries_4_specialOp_string;
  `endif


  assign _zz_stage_availROBMask_1 = (tail_0 + _zz_stage_availROBMask_2);
  assign _zz_stage_availROBMask_2 = {3'd0, dispatchNum};
  assign _zz_stage_availROBMask_4 = (tail_1 + _zz_stage_availROBMask_5);
  assign _zz_stage_availROBMask_5 = {3'd0, dispatchNum};
  assign _zz_tail_0 = (tail_0 + _zz_tail_0_1);
  assign _zz_tail_0_1 = {3'd0, dispatchNum};
  assign _zz_tail_1_1 = 1'b1;
  assign _zz_tail_1 = {4'd0, _zz_tail_1_1};
  assign _zz_tail_1_2 = (tail_1 + _zz_tail_1_3);
  assign _zz_tail_1_3 = {3'd0, dispatchNum};
  assign _zz_head_0 = (head_0 + _zz_head_0_1);
  assign _zz_head_0_1 = {3'd0, retireNum};
  assign _zz_head_1 = (head_1 + _zz_head_1_1);
  assign _zz_head_1_1 = {3'd0, retireNum};
  assign _zz_noPPRDMaskMid_1_0 = {noPPRDMaskMid_0_1,noPPRDMaskMid_0_0};
  assign _zz_freePRFIdxMid_1_0 = {noPPRDMaskMid_0_1,noPPRDMaskMid_0_0};
  assign _zz_noPPRDMaskMid_1_1 = {noPPRDMaskMid_0_1,noPPRDMaskMid_0_0};
  assign _zz_freePRFIdxMid_1_1 = {noPPRDMaskMid_0_1,noPPRDMaskMid_0_0};
  assign _zz_dispatchNum_1 = {io_dispatch_allowMask[1],io_dispatch_allowMask[0]};
  assign _zz_retireNum_1 = {retireMask[1],retireMask[0]};
  assign _zz_stage_freePRFNum_2 = {_zz_stage_freePRFNum[1],_zz_stage_freePRFNum[0]};
  always @(*) begin
    case(head_0)
      5'b00000 : begin
        _zz__zz_retirePC_0 = rob_0_pc;
        _zz__zz_noPPRDMask = rob_0_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_0_specialOp;
        _zz__zz_retireMask = rob_0_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_0_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_0_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_0_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_0_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_0_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_0_valid;
        _zz_stage_retireARAT_0_ard = rob_0_ard;
        _zz_stage_retireARAT_0_prd = rob_0_prd;
        _zz_retireTargetPC_0 = rob_0_branchResult_targetPC;
      end
      5'b00001 : begin
        _zz__zz_retirePC_0 = rob_1_pc;
        _zz__zz_noPPRDMask = rob_1_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_1_specialOp;
        _zz__zz_retireMask = rob_1_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_1_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_1_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_1_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_1_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_1_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_1_valid;
        _zz_stage_retireARAT_0_ard = rob_1_ard;
        _zz_stage_retireARAT_0_prd = rob_1_prd;
        _zz_retireTargetPC_0 = rob_1_branchResult_targetPC;
      end
      5'b00010 : begin
        _zz__zz_retirePC_0 = rob_2_pc;
        _zz__zz_noPPRDMask = rob_2_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_2_specialOp;
        _zz__zz_retireMask = rob_2_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_2_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_2_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_2_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_2_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_2_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_2_valid;
        _zz_stage_retireARAT_0_ard = rob_2_ard;
        _zz_stage_retireARAT_0_prd = rob_2_prd;
        _zz_retireTargetPC_0 = rob_2_branchResult_targetPC;
      end
      5'b00011 : begin
        _zz__zz_retirePC_0 = rob_3_pc;
        _zz__zz_noPPRDMask = rob_3_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_3_specialOp;
        _zz__zz_retireMask = rob_3_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_3_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_3_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_3_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_3_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_3_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_3_valid;
        _zz_stage_retireARAT_0_ard = rob_3_ard;
        _zz_stage_retireARAT_0_prd = rob_3_prd;
        _zz_retireTargetPC_0 = rob_3_branchResult_targetPC;
      end
      5'b00100 : begin
        _zz__zz_retirePC_0 = rob_4_pc;
        _zz__zz_noPPRDMask = rob_4_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_4_specialOp;
        _zz__zz_retireMask = rob_4_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_4_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_4_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_4_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_4_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_4_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_4_valid;
        _zz_stage_retireARAT_0_ard = rob_4_ard;
        _zz_stage_retireARAT_0_prd = rob_4_prd;
        _zz_retireTargetPC_0 = rob_4_branchResult_targetPC;
      end
      5'b00101 : begin
        _zz__zz_retirePC_0 = rob_5_pc;
        _zz__zz_noPPRDMask = rob_5_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_5_specialOp;
        _zz__zz_retireMask = rob_5_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_5_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_5_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_5_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_5_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_5_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_5_valid;
        _zz_stage_retireARAT_0_ard = rob_5_ard;
        _zz_stage_retireARAT_0_prd = rob_5_prd;
        _zz_retireTargetPC_0 = rob_5_branchResult_targetPC;
      end
      5'b00110 : begin
        _zz__zz_retirePC_0 = rob_6_pc;
        _zz__zz_noPPRDMask = rob_6_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_6_specialOp;
        _zz__zz_retireMask = rob_6_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_6_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_6_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_6_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_6_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_6_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_6_valid;
        _zz_stage_retireARAT_0_ard = rob_6_ard;
        _zz_stage_retireARAT_0_prd = rob_6_prd;
        _zz_retireTargetPC_0 = rob_6_branchResult_targetPC;
      end
      5'b00111 : begin
        _zz__zz_retirePC_0 = rob_7_pc;
        _zz__zz_noPPRDMask = rob_7_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_7_specialOp;
        _zz__zz_retireMask = rob_7_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_7_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_7_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_7_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_7_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_7_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_7_valid;
        _zz_stage_retireARAT_0_ard = rob_7_ard;
        _zz_stage_retireARAT_0_prd = rob_7_prd;
        _zz_retireTargetPC_0 = rob_7_branchResult_targetPC;
      end
      5'b01000 : begin
        _zz__zz_retirePC_0 = rob_8_pc;
        _zz__zz_noPPRDMask = rob_8_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_8_specialOp;
        _zz__zz_retireMask = rob_8_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_8_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_8_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_8_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_8_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_8_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_8_valid;
        _zz_stage_retireARAT_0_ard = rob_8_ard;
        _zz_stage_retireARAT_0_prd = rob_8_prd;
        _zz_retireTargetPC_0 = rob_8_branchResult_targetPC;
      end
      5'b01001 : begin
        _zz__zz_retirePC_0 = rob_9_pc;
        _zz__zz_noPPRDMask = rob_9_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_9_specialOp;
        _zz__zz_retireMask = rob_9_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_9_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_9_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_9_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_9_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_9_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_9_valid;
        _zz_stage_retireARAT_0_ard = rob_9_ard;
        _zz_stage_retireARAT_0_prd = rob_9_prd;
        _zz_retireTargetPC_0 = rob_9_branchResult_targetPC;
      end
      5'b01010 : begin
        _zz__zz_retirePC_0 = rob_10_pc;
        _zz__zz_noPPRDMask = rob_10_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_10_specialOp;
        _zz__zz_retireMask = rob_10_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_10_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_10_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_10_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_10_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_10_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_10_valid;
        _zz_stage_retireARAT_0_ard = rob_10_ard;
        _zz_stage_retireARAT_0_prd = rob_10_prd;
        _zz_retireTargetPC_0 = rob_10_branchResult_targetPC;
      end
      5'b01011 : begin
        _zz__zz_retirePC_0 = rob_11_pc;
        _zz__zz_noPPRDMask = rob_11_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_11_specialOp;
        _zz__zz_retireMask = rob_11_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_11_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_11_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_11_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_11_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_11_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_11_valid;
        _zz_stage_retireARAT_0_ard = rob_11_ard;
        _zz_stage_retireARAT_0_prd = rob_11_prd;
        _zz_retireTargetPC_0 = rob_11_branchResult_targetPC;
      end
      5'b01100 : begin
        _zz__zz_retirePC_0 = rob_12_pc;
        _zz__zz_noPPRDMask = rob_12_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_12_specialOp;
        _zz__zz_retireMask = rob_12_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_12_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_12_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_12_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_12_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_12_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_12_valid;
        _zz_stage_retireARAT_0_ard = rob_12_ard;
        _zz_stage_retireARAT_0_prd = rob_12_prd;
        _zz_retireTargetPC_0 = rob_12_branchResult_targetPC;
      end
      5'b01101 : begin
        _zz__zz_retirePC_0 = rob_13_pc;
        _zz__zz_noPPRDMask = rob_13_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_13_specialOp;
        _zz__zz_retireMask = rob_13_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_13_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_13_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_13_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_13_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_13_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_13_valid;
        _zz_stage_retireARAT_0_ard = rob_13_ard;
        _zz_stage_retireARAT_0_prd = rob_13_prd;
        _zz_retireTargetPC_0 = rob_13_branchResult_targetPC;
      end
      5'b01110 : begin
        _zz__zz_retirePC_0 = rob_14_pc;
        _zz__zz_noPPRDMask = rob_14_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_14_specialOp;
        _zz__zz_retireMask = rob_14_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_14_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_14_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_14_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_14_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_14_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_14_valid;
        _zz_stage_retireARAT_0_ard = rob_14_ard;
        _zz_stage_retireARAT_0_prd = rob_14_prd;
        _zz_retireTargetPC_0 = rob_14_branchResult_targetPC;
      end
      5'b01111 : begin
        _zz__zz_retirePC_0 = rob_15_pc;
        _zz__zz_noPPRDMask = rob_15_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_15_specialOp;
        _zz__zz_retireMask = rob_15_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_15_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_15_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_15_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_15_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_15_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_15_valid;
        _zz_stage_retireARAT_0_ard = rob_15_ard;
        _zz_stage_retireARAT_0_prd = rob_15_prd;
        _zz_retireTargetPC_0 = rob_15_branchResult_targetPC;
      end
      5'b10000 : begin
        _zz__zz_retirePC_0 = rob_16_pc;
        _zz__zz_noPPRDMask = rob_16_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_16_specialOp;
        _zz__zz_retireMask = rob_16_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_16_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_16_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_16_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_16_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_16_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_16_valid;
        _zz_stage_retireARAT_0_ard = rob_16_ard;
        _zz_stage_retireARAT_0_prd = rob_16_prd;
        _zz_retireTargetPC_0 = rob_16_branchResult_targetPC;
      end
      5'b10001 : begin
        _zz__zz_retirePC_0 = rob_17_pc;
        _zz__zz_noPPRDMask = rob_17_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_17_specialOp;
        _zz__zz_retireMask = rob_17_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_17_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_17_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_17_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_17_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_17_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_17_valid;
        _zz_stage_retireARAT_0_ard = rob_17_ard;
        _zz_stage_retireARAT_0_prd = rob_17_prd;
        _zz_retireTargetPC_0 = rob_17_branchResult_targetPC;
      end
      5'b10010 : begin
        _zz__zz_retirePC_0 = rob_18_pc;
        _zz__zz_noPPRDMask = rob_18_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_18_specialOp;
        _zz__zz_retireMask = rob_18_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_18_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_18_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_18_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_18_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_18_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_18_valid;
        _zz_stage_retireARAT_0_ard = rob_18_ard;
        _zz_stage_retireARAT_0_prd = rob_18_prd;
        _zz_retireTargetPC_0 = rob_18_branchResult_targetPC;
      end
      5'b10011 : begin
        _zz__zz_retirePC_0 = rob_19_pc;
        _zz__zz_noPPRDMask = rob_19_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_19_specialOp;
        _zz__zz_retireMask = rob_19_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_19_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_19_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_19_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_19_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_19_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_19_valid;
        _zz_stage_retireARAT_0_ard = rob_19_ard;
        _zz_stage_retireARAT_0_prd = rob_19_prd;
        _zz_retireTargetPC_0 = rob_19_branchResult_targetPC;
      end
      5'b10100 : begin
        _zz__zz_retirePC_0 = rob_20_pc;
        _zz__zz_noPPRDMask = rob_20_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_20_specialOp;
        _zz__zz_retireMask = rob_20_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_20_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_20_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_20_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_20_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_20_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_20_valid;
        _zz_stage_retireARAT_0_ard = rob_20_ard;
        _zz_stage_retireARAT_0_prd = rob_20_prd;
        _zz_retireTargetPC_0 = rob_20_branchResult_targetPC;
      end
      5'b10101 : begin
        _zz__zz_retirePC_0 = rob_21_pc;
        _zz__zz_noPPRDMask = rob_21_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_21_specialOp;
        _zz__zz_retireMask = rob_21_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_21_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_21_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_21_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_21_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_21_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_21_valid;
        _zz_stage_retireARAT_0_ard = rob_21_ard;
        _zz_stage_retireARAT_0_prd = rob_21_prd;
        _zz_retireTargetPC_0 = rob_21_branchResult_targetPC;
      end
      5'b10110 : begin
        _zz__zz_retirePC_0 = rob_22_pc;
        _zz__zz_noPPRDMask = rob_22_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_22_specialOp;
        _zz__zz_retireMask = rob_22_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_22_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_22_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_22_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_22_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_22_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_22_valid;
        _zz_stage_retireARAT_0_ard = rob_22_ard;
        _zz_stage_retireARAT_0_prd = rob_22_prd;
        _zz_retireTargetPC_0 = rob_22_branchResult_targetPC;
      end
      5'b10111 : begin
        _zz__zz_retirePC_0 = rob_23_pc;
        _zz__zz_noPPRDMask = rob_23_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_23_specialOp;
        _zz__zz_retireMask = rob_23_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_23_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_23_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_23_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_23_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_23_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_23_valid;
        _zz_stage_retireARAT_0_ard = rob_23_ard;
        _zz_stage_retireARAT_0_prd = rob_23_prd;
        _zz_retireTargetPC_0 = rob_23_branchResult_targetPC;
      end
      5'b11000 : begin
        _zz__zz_retirePC_0 = rob_24_pc;
        _zz__zz_noPPRDMask = rob_24_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_24_specialOp;
        _zz__zz_retireMask = rob_24_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_24_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_24_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_24_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_24_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_24_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_24_valid;
        _zz_stage_retireARAT_0_ard = rob_24_ard;
        _zz_stage_retireARAT_0_prd = rob_24_prd;
        _zz_retireTargetPC_0 = rob_24_branchResult_targetPC;
      end
      5'b11001 : begin
        _zz__zz_retirePC_0 = rob_25_pc;
        _zz__zz_noPPRDMask = rob_25_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_25_specialOp;
        _zz__zz_retireMask = rob_25_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_25_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_25_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_25_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_25_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_25_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_25_valid;
        _zz_stage_retireARAT_0_ard = rob_25_ard;
        _zz_stage_retireARAT_0_prd = rob_25_prd;
        _zz_retireTargetPC_0 = rob_25_branchResult_targetPC;
      end
      5'b11010 : begin
        _zz__zz_retirePC_0 = rob_26_pc;
        _zz__zz_noPPRDMask = rob_26_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_26_specialOp;
        _zz__zz_retireMask = rob_26_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_26_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_26_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_26_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_26_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_26_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_26_valid;
        _zz_stage_retireARAT_0_ard = rob_26_ard;
        _zz_stage_retireARAT_0_prd = rob_26_prd;
        _zz_retireTargetPC_0 = rob_26_branchResult_targetPC;
      end
      5'b11011 : begin
        _zz__zz_retirePC_0 = rob_27_pc;
        _zz__zz_noPPRDMask = rob_27_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_27_specialOp;
        _zz__zz_retireMask = rob_27_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_27_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_27_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_27_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_27_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_27_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_27_valid;
        _zz_stage_retireARAT_0_ard = rob_27_ard;
        _zz_stage_retireARAT_0_prd = rob_27_prd;
        _zz_retireTargetPC_0 = rob_27_branchResult_targetPC;
      end
      5'b11100 : begin
        _zz__zz_retirePC_0 = rob_28_pc;
        _zz__zz_noPPRDMask = rob_28_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_28_specialOp;
        _zz__zz_retireMask = rob_28_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_28_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_28_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_28_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_28_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_28_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_28_valid;
        _zz_stage_retireARAT_0_ard = rob_28_ard;
        _zz_stage_retireARAT_0_prd = rob_28_prd;
        _zz_retireTargetPC_0 = rob_28_branchResult_targetPC;
      end
      5'b11101 : begin
        _zz__zz_retirePC_0 = rob_29_pc;
        _zz__zz_noPPRDMask = rob_29_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_29_specialOp;
        _zz__zz_retireMask = rob_29_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_29_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_29_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_29_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_29_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_29_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_29_valid;
        _zz_stage_retireARAT_0_ard = rob_29_ard;
        _zz_stage_retireARAT_0_prd = rob_29_prd;
        _zz_retireTargetPC_0 = rob_29_branchResult_targetPC;
      end
      5'b11110 : begin
        _zz__zz_retirePC_0 = rob_30_pc;
        _zz__zz_noPPRDMask = rob_30_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_30_specialOp;
        _zz__zz_retireMask = rob_30_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_30_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_30_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_30_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_30_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_30_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_30_valid;
        _zz_stage_retireARAT_0_ard = rob_30_ard;
        _zz_stage_retireARAT_0_prd = rob_30_prd;
        _zz_retireTargetPC_0 = rob_30_branchResult_targetPC;
      end
      default : begin
        _zz__zz_retirePC_0 = rob_31_pc;
        _zz__zz_noPPRDMask = rob_31_pprd;
        _zz__zz_stage_updateBPU_0_isJumpInst = rob_31_specialOp;
        _zz__zz_retireMask = rob_31_isComplete;
        _zz__zz_stage_updateBPU_0_taken = rob_31_branchResult_branchResult;
        _zz__zz_stage_updateBPU_0_predictFail = rob_31_branchResult_predictFail;
        _zz__zz_retireMask_1 = rob_31_exceptionInfo_exception;
        _zz__zz_normalExceptionMask = rob_31_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_1 = rob_31_exceptionInfo_eSubCode;
        _zz__zz_retireMask_2 = rob_31_valid;
        _zz_stage_retireARAT_0_ard = rob_31_ard;
        _zz_stage_retireARAT_0_prd = rob_31_prd;
        _zz_retireTargetPC_0 = rob_31_branchResult_targetPC;
      end
    endcase
  end

  always @(*) begin
    case(_zz_dispatchNum_1)
      2'b00 : _zz_dispatchNum = 2'b00;
      2'b01 : _zz_dispatchNum = 2'b01;
      2'b10 : _zz_dispatchNum = 2'b01;
      default : _zz_dispatchNum = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_retireNum_1)
      2'b00 : _zz_retireNum = 2'b00;
      2'b01 : _zz_retireNum = 2'b01;
      2'b10 : _zz_retireNum = 2'b01;
      default : _zz_retireNum = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_stage_availROBMask_1)
      5'b00000 : _zz_stage_availROBMask = rob_0_valid;
      5'b00001 : _zz_stage_availROBMask = rob_1_valid;
      5'b00010 : _zz_stage_availROBMask = rob_2_valid;
      5'b00011 : _zz_stage_availROBMask = rob_3_valid;
      5'b00100 : _zz_stage_availROBMask = rob_4_valid;
      5'b00101 : _zz_stage_availROBMask = rob_5_valid;
      5'b00110 : _zz_stage_availROBMask = rob_6_valid;
      5'b00111 : _zz_stage_availROBMask = rob_7_valid;
      5'b01000 : _zz_stage_availROBMask = rob_8_valid;
      5'b01001 : _zz_stage_availROBMask = rob_9_valid;
      5'b01010 : _zz_stage_availROBMask = rob_10_valid;
      5'b01011 : _zz_stage_availROBMask = rob_11_valid;
      5'b01100 : _zz_stage_availROBMask = rob_12_valid;
      5'b01101 : _zz_stage_availROBMask = rob_13_valid;
      5'b01110 : _zz_stage_availROBMask = rob_14_valid;
      5'b01111 : _zz_stage_availROBMask = rob_15_valid;
      5'b10000 : _zz_stage_availROBMask = rob_16_valid;
      5'b10001 : _zz_stage_availROBMask = rob_17_valid;
      5'b10010 : _zz_stage_availROBMask = rob_18_valid;
      5'b10011 : _zz_stage_availROBMask = rob_19_valid;
      5'b10100 : _zz_stage_availROBMask = rob_20_valid;
      5'b10101 : _zz_stage_availROBMask = rob_21_valid;
      5'b10110 : _zz_stage_availROBMask = rob_22_valid;
      5'b10111 : _zz_stage_availROBMask = rob_23_valid;
      5'b11000 : _zz_stage_availROBMask = rob_24_valid;
      5'b11001 : _zz_stage_availROBMask = rob_25_valid;
      5'b11010 : _zz_stage_availROBMask = rob_26_valid;
      5'b11011 : _zz_stage_availROBMask = rob_27_valid;
      5'b11100 : _zz_stage_availROBMask = rob_28_valid;
      5'b11101 : _zz_stage_availROBMask = rob_29_valid;
      5'b11110 : _zz_stage_availROBMask = rob_30_valid;
      default : _zz_stage_availROBMask = rob_31_valid;
    endcase
  end

  always @(*) begin
    case(_zz_stage_availROBMask_4)
      5'b00000 : _zz_stage_availROBMask_3 = rob_0_valid;
      5'b00001 : _zz_stage_availROBMask_3 = rob_1_valid;
      5'b00010 : _zz_stage_availROBMask_3 = rob_2_valid;
      5'b00011 : _zz_stage_availROBMask_3 = rob_3_valid;
      5'b00100 : _zz_stage_availROBMask_3 = rob_4_valid;
      5'b00101 : _zz_stage_availROBMask_3 = rob_5_valid;
      5'b00110 : _zz_stage_availROBMask_3 = rob_6_valid;
      5'b00111 : _zz_stage_availROBMask_3 = rob_7_valid;
      5'b01000 : _zz_stage_availROBMask_3 = rob_8_valid;
      5'b01001 : _zz_stage_availROBMask_3 = rob_9_valid;
      5'b01010 : _zz_stage_availROBMask_3 = rob_10_valid;
      5'b01011 : _zz_stage_availROBMask_3 = rob_11_valid;
      5'b01100 : _zz_stage_availROBMask_3 = rob_12_valid;
      5'b01101 : _zz_stage_availROBMask_3 = rob_13_valid;
      5'b01110 : _zz_stage_availROBMask_3 = rob_14_valid;
      5'b01111 : _zz_stage_availROBMask_3 = rob_15_valid;
      5'b10000 : _zz_stage_availROBMask_3 = rob_16_valid;
      5'b10001 : _zz_stage_availROBMask_3 = rob_17_valid;
      5'b10010 : _zz_stage_availROBMask_3 = rob_18_valid;
      5'b10011 : _zz_stage_availROBMask_3 = rob_19_valid;
      5'b10100 : _zz_stage_availROBMask_3 = rob_20_valid;
      5'b10101 : _zz_stage_availROBMask_3 = rob_21_valid;
      5'b10110 : _zz_stage_availROBMask_3 = rob_22_valid;
      5'b10111 : _zz_stage_availROBMask_3 = rob_23_valid;
      5'b11000 : _zz_stage_availROBMask_3 = rob_24_valid;
      5'b11001 : _zz_stage_availROBMask_3 = rob_25_valid;
      5'b11010 : _zz_stage_availROBMask_3 = rob_26_valid;
      5'b11011 : _zz_stage_availROBMask_3 = rob_27_valid;
      5'b11100 : _zz_stage_availROBMask_3 = rob_28_valid;
      5'b11101 : _zz_stage_availROBMask_3 = rob_29_valid;
      5'b11110 : _zz_stage_availROBMask_3 = rob_30_valid;
      default : _zz_stage_availROBMask_3 = rob_31_valid;
    endcase
  end

  always @(*) begin
    case(head_1)
      5'b00000 : begin
        _zz__zz_retirePC_1 = rob_0_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_0_specialOp;
        _zz__zz_retireMask_3 = rob_0_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_0_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_0_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_0_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_0_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_0_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_0_valid;
        _zz_stage_retireARAT_1_ard = rob_0_ard;
        _zz_stage_retireARAT_1_prd = rob_0_prd;
        _zz_noPPRDMask_1 = rob_0_pprd;
        _zz_retireTargetPC_1 = rob_0_branchResult_targetPC;
      end
      5'b00001 : begin
        _zz__zz_retirePC_1 = rob_1_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_1_specialOp;
        _zz__zz_retireMask_3 = rob_1_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_1_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_1_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_1_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_1_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_1_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_1_valid;
        _zz_stage_retireARAT_1_ard = rob_1_ard;
        _zz_stage_retireARAT_1_prd = rob_1_prd;
        _zz_noPPRDMask_1 = rob_1_pprd;
        _zz_retireTargetPC_1 = rob_1_branchResult_targetPC;
      end
      5'b00010 : begin
        _zz__zz_retirePC_1 = rob_2_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_2_specialOp;
        _zz__zz_retireMask_3 = rob_2_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_2_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_2_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_2_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_2_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_2_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_2_valid;
        _zz_stage_retireARAT_1_ard = rob_2_ard;
        _zz_stage_retireARAT_1_prd = rob_2_prd;
        _zz_noPPRDMask_1 = rob_2_pprd;
        _zz_retireTargetPC_1 = rob_2_branchResult_targetPC;
      end
      5'b00011 : begin
        _zz__zz_retirePC_1 = rob_3_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_3_specialOp;
        _zz__zz_retireMask_3 = rob_3_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_3_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_3_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_3_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_3_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_3_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_3_valid;
        _zz_stage_retireARAT_1_ard = rob_3_ard;
        _zz_stage_retireARAT_1_prd = rob_3_prd;
        _zz_noPPRDMask_1 = rob_3_pprd;
        _zz_retireTargetPC_1 = rob_3_branchResult_targetPC;
      end
      5'b00100 : begin
        _zz__zz_retirePC_1 = rob_4_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_4_specialOp;
        _zz__zz_retireMask_3 = rob_4_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_4_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_4_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_4_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_4_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_4_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_4_valid;
        _zz_stage_retireARAT_1_ard = rob_4_ard;
        _zz_stage_retireARAT_1_prd = rob_4_prd;
        _zz_noPPRDMask_1 = rob_4_pprd;
        _zz_retireTargetPC_1 = rob_4_branchResult_targetPC;
      end
      5'b00101 : begin
        _zz__zz_retirePC_1 = rob_5_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_5_specialOp;
        _zz__zz_retireMask_3 = rob_5_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_5_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_5_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_5_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_5_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_5_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_5_valid;
        _zz_stage_retireARAT_1_ard = rob_5_ard;
        _zz_stage_retireARAT_1_prd = rob_5_prd;
        _zz_noPPRDMask_1 = rob_5_pprd;
        _zz_retireTargetPC_1 = rob_5_branchResult_targetPC;
      end
      5'b00110 : begin
        _zz__zz_retirePC_1 = rob_6_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_6_specialOp;
        _zz__zz_retireMask_3 = rob_6_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_6_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_6_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_6_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_6_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_6_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_6_valid;
        _zz_stage_retireARAT_1_ard = rob_6_ard;
        _zz_stage_retireARAT_1_prd = rob_6_prd;
        _zz_noPPRDMask_1 = rob_6_pprd;
        _zz_retireTargetPC_1 = rob_6_branchResult_targetPC;
      end
      5'b00111 : begin
        _zz__zz_retirePC_1 = rob_7_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_7_specialOp;
        _zz__zz_retireMask_3 = rob_7_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_7_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_7_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_7_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_7_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_7_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_7_valid;
        _zz_stage_retireARAT_1_ard = rob_7_ard;
        _zz_stage_retireARAT_1_prd = rob_7_prd;
        _zz_noPPRDMask_1 = rob_7_pprd;
        _zz_retireTargetPC_1 = rob_7_branchResult_targetPC;
      end
      5'b01000 : begin
        _zz__zz_retirePC_1 = rob_8_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_8_specialOp;
        _zz__zz_retireMask_3 = rob_8_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_8_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_8_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_8_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_8_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_8_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_8_valid;
        _zz_stage_retireARAT_1_ard = rob_8_ard;
        _zz_stage_retireARAT_1_prd = rob_8_prd;
        _zz_noPPRDMask_1 = rob_8_pprd;
        _zz_retireTargetPC_1 = rob_8_branchResult_targetPC;
      end
      5'b01001 : begin
        _zz__zz_retirePC_1 = rob_9_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_9_specialOp;
        _zz__zz_retireMask_3 = rob_9_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_9_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_9_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_9_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_9_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_9_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_9_valid;
        _zz_stage_retireARAT_1_ard = rob_9_ard;
        _zz_stage_retireARAT_1_prd = rob_9_prd;
        _zz_noPPRDMask_1 = rob_9_pprd;
        _zz_retireTargetPC_1 = rob_9_branchResult_targetPC;
      end
      5'b01010 : begin
        _zz__zz_retirePC_1 = rob_10_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_10_specialOp;
        _zz__zz_retireMask_3 = rob_10_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_10_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_10_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_10_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_10_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_10_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_10_valid;
        _zz_stage_retireARAT_1_ard = rob_10_ard;
        _zz_stage_retireARAT_1_prd = rob_10_prd;
        _zz_noPPRDMask_1 = rob_10_pprd;
        _zz_retireTargetPC_1 = rob_10_branchResult_targetPC;
      end
      5'b01011 : begin
        _zz__zz_retirePC_1 = rob_11_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_11_specialOp;
        _zz__zz_retireMask_3 = rob_11_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_11_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_11_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_11_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_11_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_11_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_11_valid;
        _zz_stage_retireARAT_1_ard = rob_11_ard;
        _zz_stage_retireARAT_1_prd = rob_11_prd;
        _zz_noPPRDMask_1 = rob_11_pprd;
        _zz_retireTargetPC_1 = rob_11_branchResult_targetPC;
      end
      5'b01100 : begin
        _zz__zz_retirePC_1 = rob_12_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_12_specialOp;
        _zz__zz_retireMask_3 = rob_12_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_12_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_12_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_12_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_12_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_12_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_12_valid;
        _zz_stage_retireARAT_1_ard = rob_12_ard;
        _zz_stage_retireARAT_1_prd = rob_12_prd;
        _zz_noPPRDMask_1 = rob_12_pprd;
        _zz_retireTargetPC_1 = rob_12_branchResult_targetPC;
      end
      5'b01101 : begin
        _zz__zz_retirePC_1 = rob_13_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_13_specialOp;
        _zz__zz_retireMask_3 = rob_13_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_13_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_13_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_13_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_13_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_13_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_13_valid;
        _zz_stage_retireARAT_1_ard = rob_13_ard;
        _zz_stage_retireARAT_1_prd = rob_13_prd;
        _zz_noPPRDMask_1 = rob_13_pprd;
        _zz_retireTargetPC_1 = rob_13_branchResult_targetPC;
      end
      5'b01110 : begin
        _zz__zz_retirePC_1 = rob_14_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_14_specialOp;
        _zz__zz_retireMask_3 = rob_14_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_14_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_14_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_14_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_14_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_14_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_14_valid;
        _zz_stage_retireARAT_1_ard = rob_14_ard;
        _zz_stage_retireARAT_1_prd = rob_14_prd;
        _zz_noPPRDMask_1 = rob_14_pprd;
        _zz_retireTargetPC_1 = rob_14_branchResult_targetPC;
      end
      5'b01111 : begin
        _zz__zz_retirePC_1 = rob_15_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_15_specialOp;
        _zz__zz_retireMask_3 = rob_15_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_15_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_15_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_15_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_15_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_15_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_15_valid;
        _zz_stage_retireARAT_1_ard = rob_15_ard;
        _zz_stage_retireARAT_1_prd = rob_15_prd;
        _zz_noPPRDMask_1 = rob_15_pprd;
        _zz_retireTargetPC_1 = rob_15_branchResult_targetPC;
      end
      5'b10000 : begin
        _zz__zz_retirePC_1 = rob_16_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_16_specialOp;
        _zz__zz_retireMask_3 = rob_16_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_16_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_16_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_16_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_16_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_16_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_16_valid;
        _zz_stage_retireARAT_1_ard = rob_16_ard;
        _zz_stage_retireARAT_1_prd = rob_16_prd;
        _zz_noPPRDMask_1 = rob_16_pprd;
        _zz_retireTargetPC_1 = rob_16_branchResult_targetPC;
      end
      5'b10001 : begin
        _zz__zz_retirePC_1 = rob_17_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_17_specialOp;
        _zz__zz_retireMask_3 = rob_17_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_17_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_17_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_17_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_17_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_17_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_17_valid;
        _zz_stage_retireARAT_1_ard = rob_17_ard;
        _zz_stage_retireARAT_1_prd = rob_17_prd;
        _zz_noPPRDMask_1 = rob_17_pprd;
        _zz_retireTargetPC_1 = rob_17_branchResult_targetPC;
      end
      5'b10010 : begin
        _zz__zz_retirePC_1 = rob_18_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_18_specialOp;
        _zz__zz_retireMask_3 = rob_18_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_18_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_18_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_18_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_18_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_18_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_18_valid;
        _zz_stage_retireARAT_1_ard = rob_18_ard;
        _zz_stage_retireARAT_1_prd = rob_18_prd;
        _zz_noPPRDMask_1 = rob_18_pprd;
        _zz_retireTargetPC_1 = rob_18_branchResult_targetPC;
      end
      5'b10011 : begin
        _zz__zz_retirePC_1 = rob_19_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_19_specialOp;
        _zz__zz_retireMask_3 = rob_19_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_19_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_19_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_19_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_19_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_19_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_19_valid;
        _zz_stage_retireARAT_1_ard = rob_19_ard;
        _zz_stage_retireARAT_1_prd = rob_19_prd;
        _zz_noPPRDMask_1 = rob_19_pprd;
        _zz_retireTargetPC_1 = rob_19_branchResult_targetPC;
      end
      5'b10100 : begin
        _zz__zz_retirePC_1 = rob_20_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_20_specialOp;
        _zz__zz_retireMask_3 = rob_20_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_20_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_20_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_20_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_20_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_20_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_20_valid;
        _zz_stage_retireARAT_1_ard = rob_20_ard;
        _zz_stage_retireARAT_1_prd = rob_20_prd;
        _zz_noPPRDMask_1 = rob_20_pprd;
        _zz_retireTargetPC_1 = rob_20_branchResult_targetPC;
      end
      5'b10101 : begin
        _zz__zz_retirePC_1 = rob_21_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_21_specialOp;
        _zz__zz_retireMask_3 = rob_21_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_21_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_21_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_21_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_21_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_21_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_21_valid;
        _zz_stage_retireARAT_1_ard = rob_21_ard;
        _zz_stage_retireARAT_1_prd = rob_21_prd;
        _zz_noPPRDMask_1 = rob_21_pprd;
        _zz_retireTargetPC_1 = rob_21_branchResult_targetPC;
      end
      5'b10110 : begin
        _zz__zz_retirePC_1 = rob_22_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_22_specialOp;
        _zz__zz_retireMask_3 = rob_22_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_22_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_22_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_22_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_22_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_22_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_22_valid;
        _zz_stage_retireARAT_1_ard = rob_22_ard;
        _zz_stage_retireARAT_1_prd = rob_22_prd;
        _zz_noPPRDMask_1 = rob_22_pprd;
        _zz_retireTargetPC_1 = rob_22_branchResult_targetPC;
      end
      5'b10111 : begin
        _zz__zz_retirePC_1 = rob_23_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_23_specialOp;
        _zz__zz_retireMask_3 = rob_23_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_23_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_23_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_23_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_23_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_23_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_23_valid;
        _zz_stage_retireARAT_1_ard = rob_23_ard;
        _zz_stage_retireARAT_1_prd = rob_23_prd;
        _zz_noPPRDMask_1 = rob_23_pprd;
        _zz_retireTargetPC_1 = rob_23_branchResult_targetPC;
      end
      5'b11000 : begin
        _zz__zz_retirePC_1 = rob_24_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_24_specialOp;
        _zz__zz_retireMask_3 = rob_24_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_24_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_24_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_24_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_24_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_24_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_24_valid;
        _zz_stage_retireARAT_1_ard = rob_24_ard;
        _zz_stage_retireARAT_1_prd = rob_24_prd;
        _zz_noPPRDMask_1 = rob_24_pprd;
        _zz_retireTargetPC_1 = rob_24_branchResult_targetPC;
      end
      5'b11001 : begin
        _zz__zz_retirePC_1 = rob_25_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_25_specialOp;
        _zz__zz_retireMask_3 = rob_25_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_25_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_25_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_25_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_25_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_25_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_25_valid;
        _zz_stage_retireARAT_1_ard = rob_25_ard;
        _zz_stage_retireARAT_1_prd = rob_25_prd;
        _zz_noPPRDMask_1 = rob_25_pprd;
        _zz_retireTargetPC_1 = rob_25_branchResult_targetPC;
      end
      5'b11010 : begin
        _zz__zz_retirePC_1 = rob_26_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_26_specialOp;
        _zz__zz_retireMask_3 = rob_26_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_26_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_26_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_26_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_26_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_26_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_26_valid;
        _zz_stage_retireARAT_1_ard = rob_26_ard;
        _zz_stage_retireARAT_1_prd = rob_26_prd;
        _zz_noPPRDMask_1 = rob_26_pprd;
        _zz_retireTargetPC_1 = rob_26_branchResult_targetPC;
      end
      5'b11011 : begin
        _zz__zz_retirePC_1 = rob_27_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_27_specialOp;
        _zz__zz_retireMask_3 = rob_27_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_27_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_27_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_27_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_27_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_27_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_27_valid;
        _zz_stage_retireARAT_1_ard = rob_27_ard;
        _zz_stage_retireARAT_1_prd = rob_27_prd;
        _zz_noPPRDMask_1 = rob_27_pprd;
        _zz_retireTargetPC_1 = rob_27_branchResult_targetPC;
      end
      5'b11100 : begin
        _zz__zz_retirePC_1 = rob_28_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_28_specialOp;
        _zz__zz_retireMask_3 = rob_28_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_28_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_28_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_28_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_28_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_28_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_28_valid;
        _zz_stage_retireARAT_1_ard = rob_28_ard;
        _zz_stage_retireARAT_1_prd = rob_28_prd;
        _zz_noPPRDMask_1 = rob_28_pprd;
        _zz_retireTargetPC_1 = rob_28_branchResult_targetPC;
      end
      5'b11101 : begin
        _zz__zz_retirePC_1 = rob_29_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_29_specialOp;
        _zz__zz_retireMask_3 = rob_29_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_29_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_29_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_29_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_29_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_29_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_29_valid;
        _zz_stage_retireARAT_1_ard = rob_29_ard;
        _zz_stage_retireARAT_1_prd = rob_29_prd;
        _zz_noPPRDMask_1 = rob_29_pprd;
        _zz_retireTargetPC_1 = rob_29_branchResult_targetPC;
      end
      5'b11110 : begin
        _zz__zz_retirePC_1 = rob_30_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_30_specialOp;
        _zz__zz_retireMask_3 = rob_30_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_30_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_30_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_30_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_30_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_30_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_30_valid;
        _zz_stage_retireARAT_1_ard = rob_30_ard;
        _zz_stage_retireARAT_1_prd = rob_30_prd;
        _zz_noPPRDMask_1 = rob_30_pprd;
        _zz_retireTargetPC_1 = rob_30_branchResult_targetPC;
      end
      default : begin
        _zz__zz_retirePC_1 = rob_31_pc;
        _zz__zz_stage_updateBPU_1_isJumpInst = rob_31_specialOp;
        _zz__zz_retireMask_3 = rob_31_isComplete;
        _zz__zz_stage_updateBPU_1_taken = rob_31_branchResult_branchResult;
        _zz__zz_stage_updateBPU_1_predictFail = rob_31_branchResult_predictFail;
        _zz__zz_retireMask_4 = rob_31_exceptionInfo_exception;
        _zz__zz_normalExceptionMask_2 = rob_31_exceptionInfo_eCode;
        _zz__zz_normalExceptionMask_3 = rob_31_exceptionInfo_eSubCode;
        _zz__zz_retireMask_5 = rob_31_valid;
        _zz_stage_retireARAT_1_ard = rob_31_ard;
        _zz_stage_retireARAT_1_prd = rob_31_prd;
        _zz_noPPRDMask_1 = rob_31_pprd;
        _zz_retireTargetPC_1 = rob_31_branchResult_targetPC;
      end
    endcase
  end

  always @(*) begin
    case(_zz_io_commitROBEntries_0_pc)
      5'b00000 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_0_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_0_pc;
        _zz_io_commitROBEntries_0_ard = rob_0_ard;
        _zz_io_commitROBEntries_0_prd = rob_0_prd;
        _zz_io_commitROBEntries_0_pprd = rob_0_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_0_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_0_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_0_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_0_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_0_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_0_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_0_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_0_valid;
      end
      5'b00001 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_1_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_1_pc;
        _zz_io_commitROBEntries_0_ard = rob_1_ard;
        _zz_io_commitROBEntries_0_prd = rob_1_prd;
        _zz_io_commitROBEntries_0_pprd = rob_1_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_1_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_1_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_1_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_1_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_1_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_1_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_1_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_1_valid;
      end
      5'b00010 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_2_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_2_pc;
        _zz_io_commitROBEntries_0_ard = rob_2_ard;
        _zz_io_commitROBEntries_0_prd = rob_2_prd;
        _zz_io_commitROBEntries_0_pprd = rob_2_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_2_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_2_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_2_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_2_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_2_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_2_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_2_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_2_valid;
      end
      5'b00011 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_3_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_3_pc;
        _zz_io_commitROBEntries_0_ard = rob_3_ard;
        _zz_io_commitROBEntries_0_prd = rob_3_prd;
        _zz_io_commitROBEntries_0_pprd = rob_3_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_3_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_3_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_3_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_3_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_3_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_3_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_3_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_3_valid;
      end
      5'b00100 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_4_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_4_pc;
        _zz_io_commitROBEntries_0_ard = rob_4_ard;
        _zz_io_commitROBEntries_0_prd = rob_4_prd;
        _zz_io_commitROBEntries_0_pprd = rob_4_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_4_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_4_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_4_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_4_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_4_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_4_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_4_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_4_valid;
      end
      5'b00101 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_5_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_5_pc;
        _zz_io_commitROBEntries_0_ard = rob_5_ard;
        _zz_io_commitROBEntries_0_prd = rob_5_prd;
        _zz_io_commitROBEntries_0_pprd = rob_5_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_5_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_5_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_5_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_5_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_5_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_5_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_5_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_5_valid;
      end
      5'b00110 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_6_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_6_pc;
        _zz_io_commitROBEntries_0_ard = rob_6_ard;
        _zz_io_commitROBEntries_0_prd = rob_6_prd;
        _zz_io_commitROBEntries_0_pprd = rob_6_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_6_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_6_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_6_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_6_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_6_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_6_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_6_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_6_valid;
      end
      5'b00111 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_7_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_7_pc;
        _zz_io_commitROBEntries_0_ard = rob_7_ard;
        _zz_io_commitROBEntries_0_prd = rob_7_prd;
        _zz_io_commitROBEntries_0_pprd = rob_7_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_7_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_7_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_7_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_7_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_7_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_7_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_7_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_7_valid;
      end
      5'b01000 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_8_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_8_pc;
        _zz_io_commitROBEntries_0_ard = rob_8_ard;
        _zz_io_commitROBEntries_0_prd = rob_8_prd;
        _zz_io_commitROBEntries_0_pprd = rob_8_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_8_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_8_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_8_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_8_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_8_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_8_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_8_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_8_valid;
      end
      5'b01001 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_9_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_9_pc;
        _zz_io_commitROBEntries_0_ard = rob_9_ard;
        _zz_io_commitROBEntries_0_prd = rob_9_prd;
        _zz_io_commitROBEntries_0_pprd = rob_9_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_9_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_9_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_9_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_9_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_9_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_9_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_9_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_9_valid;
      end
      5'b01010 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_10_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_10_pc;
        _zz_io_commitROBEntries_0_ard = rob_10_ard;
        _zz_io_commitROBEntries_0_prd = rob_10_prd;
        _zz_io_commitROBEntries_0_pprd = rob_10_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_10_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_10_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_10_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_10_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_10_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_10_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_10_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_10_valid;
      end
      5'b01011 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_11_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_11_pc;
        _zz_io_commitROBEntries_0_ard = rob_11_ard;
        _zz_io_commitROBEntries_0_prd = rob_11_prd;
        _zz_io_commitROBEntries_0_pprd = rob_11_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_11_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_11_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_11_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_11_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_11_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_11_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_11_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_11_valid;
      end
      5'b01100 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_12_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_12_pc;
        _zz_io_commitROBEntries_0_ard = rob_12_ard;
        _zz_io_commitROBEntries_0_prd = rob_12_prd;
        _zz_io_commitROBEntries_0_pprd = rob_12_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_12_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_12_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_12_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_12_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_12_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_12_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_12_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_12_valid;
      end
      5'b01101 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_13_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_13_pc;
        _zz_io_commitROBEntries_0_ard = rob_13_ard;
        _zz_io_commitROBEntries_0_prd = rob_13_prd;
        _zz_io_commitROBEntries_0_pprd = rob_13_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_13_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_13_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_13_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_13_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_13_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_13_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_13_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_13_valid;
      end
      5'b01110 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_14_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_14_pc;
        _zz_io_commitROBEntries_0_ard = rob_14_ard;
        _zz_io_commitROBEntries_0_prd = rob_14_prd;
        _zz_io_commitROBEntries_0_pprd = rob_14_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_14_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_14_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_14_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_14_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_14_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_14_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_14_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_14_valid;
      end
      5'b01111 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_15_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_15_pc;
        _zz_io_commitROBEntries_0_ard = rob_15_ard;
        _zz_io_commitROBEntries_0_prd = rob_15_prd;
        _zz_io_commitROBEntries_0_pprd = rob_15_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_15_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_15_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_15_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_15_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_15_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_15_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_15_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_15_valid;
      end
      5'b10000 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_16_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_16_pc;
        _zz_io_commitROBEntries_0_ard = rob_16_ard;
        _zz_io_commitROBEntries_0_prd = rob_16_prd;
        _zz_io_commitROBEntries_0_pprd = rob_16_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_16_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_16_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_16_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_16_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_16_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_16_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_16_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_16_valid;
      end
      5'b10001 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_17_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_17_pc;
        _zz_io_commitROBEntries_0_ard = rob_17_ard;
        _zz_io_commitROBEntries_0_prd = rob_17_prd;
        _zz_io_commitROBEntries_0_pprd = rob_17_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_17_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_17_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_17_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_17_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_17_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_17_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_17_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_17_valid;
      end
      5'b10010 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_18_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_18_pc;
        _zz_io_commitROBEntries_0_ard = rob_18_ard;
        _zz_io_commitROBEntries_0_prd = rob_18_prd;
        _zz_io_commitROBEntries_0_pprd = rob_18_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_18_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_18_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_18_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_18_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_18_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_18_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_18_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_18_valid;
      end
      5'b10011 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_19_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_19_pc;
        _zz_io_commitROBEntries_0_ard = rob_19_ard;
        _zz_io_commitROBEntries_0_prd = rob_19_prd;
        _zz_io_commitROBEntries_0_pprd = rob_19_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_19_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_19_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_19_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_19_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_19_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_19_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_19_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_19_valid;
      end
      5'b10100 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_20_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_20_pc;
        _zz_io_commitROBEntries_0_ard = rob_20_ard;
        _zz_io_commitROBEntries_0_prd = rob_20_prd;
        _zz_io_commitROBEntries_0_pprd = rob_20_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_20_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_20_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_20_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_20_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_20_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_20_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_20_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_20_valid;
      end
      5'b10101 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_21_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_21_pc;
        _zz_io_commitROBEntries_0_ard = rob_21_ard;
        _zz_io_commitROBEntries_0_prd = rob_21_prd;
        _zz_io_commitROBEntries_0_pprd = rob_21_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_21_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_21_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_21_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_21_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_21_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_21_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_21_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_21_valid;
      end
      5'b10110 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_22_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_22_pc;
        _zz_io_commitROBEntries_0_ard = rob_22_ard;
        _zz_io_commitROBEntries_0_prd = rob_22_prd;
        _zz_io_commitROBEntries_0_pprd = rob_22_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_22_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_22_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_22_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_22_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_22_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_22_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_22_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_22_valid;
      end
      5'b10111 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_23_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_23_pc;
        _zz_io_commitROBEntries_0_ard = rob_23_ard;
        _zz_io_commitROBEntries_0_prd = rob_23_prd;
        _zz_io_commitROBEntries_0_pprd = rob_23_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_23_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_23_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_23_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_23_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_23_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_23_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_23_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_23_valid;
      end
      5'b11000 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_24_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_24_pc;
        _zz_io_commitROBEntries_0_ard = rob_24_ard;
        _zz_io_commitROBEntries_0_prd = rob_24_prd;
        _zz_io_commitROBEntries_0_pprd = rob_24_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_24_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_24_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_24_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_24_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_24_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_24_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_24_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_24_valid;
      end
      5'b11001 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_25_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_25_pc;
        _zz_io_commitROBEntries_0_ard = rob_25_ard;
        _zz_io_commitROBEntries_0_prd = rob_25_prd;
        _zz_io_commitROBEntries_0_pprd = rob_25_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_25_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_25_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_25_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_25_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_25_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_25_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_25_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_25_valid;
      end
      5'b11010 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_26_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_26_pc;
        _zz_io_commitROBEntries_0_ard = rob_26_ard;
        _zz_io_commitROBEntries_0_prd = rob_26_prd;
        _zz_io_commitROBEntries_0_pprd = rob_26_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_26_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_26_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_26_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_26_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_26_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_26_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_26_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_26_valid;
      end
      5'b11011 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_27_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_27_pc;
        _zz_io_commitROBEntries_0_ard = rob_27_ard;
        _zz_io_commitROBEntries_0_prd = rob_27_prd;
        _zz_io_commitROBEntries_0_pprd = rob_27_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_27_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_27_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_27_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_27_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_27_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_27_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_27_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_27_valid;
      end
      5'b11100 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_28_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_28_pc;
        _zz_io_commitROBEntries_0_ard = rob_28_ard;
        _zz_io_commitROBEntries_0_prd = rob_28_prd;
        _zz_io_commitROBEntries_0_pprd = rob_28_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_28_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_28_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_28_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_28_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_28_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_28_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_28_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_28_valid;
      end
      5'b11101 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_29_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_29_pc;
        _zz_io_commitROBEntries_0_ard = rob_29_ard;
        _zz_io_commitROBEntries_0_prd = rob_29_prd;
        _zz_io_commitROBEntries_0_pprd = rob_29_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_29_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_29_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_29_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_29_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_29_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_29_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_29_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_29_valid;
      end
      5'b11110 : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_30_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_30_pc;
        _zz_io_commitROBEntries_0_ard = rob_30_ard;
        _zz_io_commitROBEntries_0_prd = rob_30_prd;
        _zz_io_commitROBEntries_0_pprd = rob_30_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_30_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_30_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_30_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_30_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_30_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_30_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_30_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_30_valid;
      end
      default : begin
        _zz__zz_io_commitROBEntries_0_specialOp = rob_31_specialOp;
        _zz_io_commitROBEntries_0_pc_1 = rob_31_pc;
        _zz_io_commitROBEntries_0_ard = rob_31_ard;
        _zz_io_commitROBEntries_0_prd = rob_31_prd;
        _zz_io_commitROBEntries_0_pprd = rob_31_pprd;
        _zz_io_commitROBEntries_0_isComplete = rob_31_isComplete;
        _zz_io_commitROBEntries_0_branchResult_targetPC = rob_31_branchResult_targetPC;
        _zz_io_commitROBEntries_0_branchResult_branchResult = rob_31_branchResult_branchResult;
        _zz_io_commitROBEntries_0_branchResult_predictFail = rob_31_branchResult_predictFail;
        _zz_io_commitROBEntries_0_exceptionInfo_exception = rob_31_exceptionInfo_exception;
        _zz_io_commitROBEntries_0_exceptionInfo_eCode = rob_31_exceptionInfo_eCode;
        _zz_io_commitROBEntries_0_exceptionInfo_eSubCode = rob_31_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_0_valid = rob_31_valid;
      end
    endcase
  end

  always @(*) begin
    case(_zz_io_commitROBEntries_1_pc)
      5'b00000 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_0_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_0_pc;
        _zz_io_commitROBEntries_1_ard = rob_0_ard;
        _zz_io_commitROBEntries_1_prd = rob_0_prd;
        _zz_io_commitROBEntries_1_pprd = rob_0_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_0_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_0_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_0_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_0_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_0_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_0_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_0_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_0_valid;
      end
      5'b00001 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_1_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_1_pc;
        _zz_io_commitROBEntries_1_ard = rob_1_ard;
        _zz_io_commitROBEntries_1_prd = rob_1_prd;
        _zz_io_commitROBEntries_1_pprd = rob_1_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_1_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_1_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_1_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_1_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_1_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_1_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_1_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_1_valid;
      end
      5'b00010 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_2_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_2_pc;
        _zz_io_commitROBEntries_1_ard = rob_2_ard;
        _zz_io_commitROBEntries_1_prd = rob_2_prd;
        _zz_io_commitROBEntries_1_pprd = rob_2_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_2_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_2_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_2_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_2_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_2_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_2_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_2_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_2_valid;
      end
      5'b00011 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_3_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_3_pc;
        _zz_io_commitROBEntries_1_ard = rob_3_ard;
        _zz_io_commitROBEntries_1_prd = rob_3_prd;
        _zz_io_commitROBEntries_1_pprd = rob_3_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_3_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_3_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_3_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_3_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_3_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_3_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_3_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_3_valid;
      end
      5'b00100 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_4_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_4_pc;
        _zz_io_commitROBEntries_1_ard = rob_4_ard;
        _zz_io_commitROBEntries_1_prd = rob_4_prd;
        _zz_io_commitROBEntries_1_pprd = rob_4_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_4_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_4_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_4_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_4_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_4_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_4_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_4_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_4_valid;
      end
      5'b00101 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_5_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_5_pc;
        _zz_io_commitROBEntries_1_ard = rob_5_ard;
        _zz_io_commitROBEntries_1_prd = rob_5_prd;
        _zz_io_commitROBEntries_1_pprd = rob_5_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_5_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_5_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_5_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_5_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_5_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_5_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_5_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_5_valid;
      end
      5'b00110 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_6_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_6_pc;
        _zz_io_commitROBEntries_1_ard = rob_6_ard;
        _zz_io_commitROBEntries_1_prd = rob_6_prd;
        _zz_io_commitROBEntries_1_pprd = rob_6_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_6_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_6_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_6_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_6_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_6_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_6_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_6_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_6_valid;
      end
      5'b00111 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_7_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_7_pc;
        _zz_io_commitROBEntries_1_ard = rob_7_ard;
        _zz_io_commitROBEntries_1_prd = rob_7_prd;
        _zz_io_commitROBEntries_1_pprd = rob_7_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_7_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_7_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_7_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_7_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_7_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_7_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_7_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_7_valid;
      end
      5'b01000 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_8_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_8_pc;
        _zz_io_commitROBEntries_1_ard = rob_8_ard;
        _zz_io_commitROBEntries_1_prd = rob_8_prd;
        _zz_io_commitROBEntries_1_pprd = rob_8_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_8_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_8_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_8_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_8_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_8_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_8_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_8_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_8_valid;
      end
      5'b01001 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_9_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_9_pc;
        _zz_io_commitROBEntries_1_ard = rob_9_ard;
        _zz_io_commitROBEntries_1_prd = rob_9_prd;
        _zz_io_commitROBEntries_1_pprd = rob_9_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_9_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_9_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_9_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_9_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_9_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_9_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_9_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_9_valid;
      end
      5'b01010 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_10_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_10_pc;
        _zz_io_commitROBEntries_1_ard = rob_10_ard;
        _zz_io_commitROBEntries_1_prd = rob_10_prd;
        _zz_io_commitROBEntries_1_pprd = rob_10_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_10_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_10_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_10_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_10_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_10_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_10_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_10_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_10_valid;
      end
      5'b01011 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_11_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_11_pc;
        _zz_io_commitROBEntries_1_ard = rob_11_ard;
        _zz_io_commitROBEntries_1_prd = rob_11_prd;
        _zz_io_commitROBEntries_1_pprd = rob_11_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_11_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_11_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_11_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_11_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_11_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_11_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_11_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_11_valid;
      end
      5'b01100 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_12_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_12_pc;
        _zz_io_commitROBEntries_1_ard = rob_12_ard;
        _zz_io_commitROBEntries_1_prd = rob_12_prd;
        _zz_io_commitROBEntries_1_pprd = rob_12_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_12_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_12_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_12_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_12_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_12_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_12_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_12_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_12_valid;
      end
      5'b01101 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_13_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_13_pc;
        _zz_io_commitROBEntries_1_ard = rob_13_ard;
        _zz_io_commitROBEntries_1_prd = rob_13_prd;
        _zz_io_commitROBEntries_1_pprd = rob_13_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_13_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_13_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_13_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_13_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_13_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_13_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_13_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_13_valid;
      end
      5'b01110 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_14_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_14_pc;
        _zz_io_commitROBEntries_1_ard = rob_14_ard;
        _zz_io_commitROBEntries_1_prd = rob_14_prd;
        _zz_io_commitROBEntries_1_pprd = rob_14_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_14_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_14_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_14_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_14_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_14_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_14_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_14_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_14_valid;
      end
      5'b01111 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_15_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_15_pc;
        _zz_io_commitROBEntries_1_ard = rob_15_ard;
        _zz_io_commitROBEntries_1_prd = rob_15_prd;
        _zz_io_commitROBEntries_1_pprd = rob_15_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_15_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_15_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_15_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_15_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_15_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_15_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_15_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_15_valid;
      end
      5'b10000 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_16_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_16_pc;
        _zz_io_commitROBEntries_1_ard = rob_16_ard;
        _zz_io_commitROBEntries_1_prd = rob_16_prd;
        _zz_io_commitROBEntries_1_pprd = rob_16_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_16_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_16_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_16_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_16_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_16_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_16_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_16_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_16_valid;
      end
      5'b10001 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_17_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_17_pc;
        _zz_io_commitROBEntries_1_ard = rob_17_ard;
        _zz_io_commitROBEntries_1_prd = rob_17_prd;
        _zz_io_commitROBEntries_1_pprd = rob_17_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_17_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_17_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_17_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_17_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_17_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_17_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_17_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_17_valid;
      end
      5'b10010 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_18_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_18_pc;
        _zz_io_commitROBEntries_1_ard = rob_18_ard;
        _zz_io_commitROBEntries_1_prd = rob_18_prd;
        _zz_io_commitROBEntries_1_pprd = rob_18_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_18_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_18_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_18_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_18_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_18_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_18_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_18_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_18_valid;
      end
      5'b10011 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_19_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_19_pc;
        _zz_io_commitROBEntries_1_ard = rob_19_ard;
        _zz_io_commitROBEntries_1_prd = rob_19_prd;
        _zz_io_commitROBEntries_1_pprd = rob_19_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_19_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_19_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_19_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_19_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_19_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_19_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_19_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_19_valid;
      end
      5'b10100 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_20_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_20_pc;
        _zz_io_commitROBEntries_1_ard = rob_20_ard;
        _zz_io_commitROBEntries_1_prd = rob_20_prd;
        _zz_io_commitROBEntries_1_pprd = rob_20_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_20_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_20_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_20_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_20_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_20_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_20_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_20_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_20_valid;
      end
      5'b10101 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_21_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_21_pc;
        _zz_io_commitROBEntries_1_ard = rob_21_ard;
        _zz_io_commitROBEntries_1_prd = rob_21_prd;
        _zz_io_commitROBEntries_1_pprd = rob_21_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_21_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_21_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_21_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_21_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_21_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_21_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_21_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_21_valid;
      end
      5'b10110 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_22_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_22_pc;
        _zz_io_commitROBEntries_1_ard = rob_22_ard;
        _zz_io_commitROBEntries_1_prd = rob_22_prd;
        _zz_io_commitROBEntries_1_pprd = rob_22_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_22_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_22_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_22_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_22_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_22_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_22_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_22_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_22_valid;
      end
      5'b10111 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_23_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_23_pc;
        _zz_io_commitROBEntries_1_ard = rob_23_ard;
        _zz_io_commitROBEntries_1_prd = rob_23_prd;
        _zz_io_commitROBEntries_1_pprd = rob_23_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_23_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_23_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_23_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_23_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_23_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_23_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_23_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_23_valid;
      end
      5'b11000 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_24_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_24_pc;
        _zz_io_commitROBEntries_1_ard = rob_24_ard;
        _zz_io_commitROBEntries_1_prd = rob_24_prd;
        _zz_io_commitROBEntries_1_pprd = rob_24_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_24_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_24_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_24_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_24_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_24_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_24_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_24_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_24_valid;
      end
      5'b11001 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_25_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_25_pc;
        _zz_io_commitROBEntries_1_ard = rob_25_ard;
        _zz_io_commitROBEntries_1_prd = rob_25_prd;
        _zz_io_commitROBEntries_1_pprd = rob_25_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_25_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_25_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_25_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_25_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_25_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_25_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_25_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_25_valid;
      end
      5'b11010 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_26_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_26_pc;
        _zz_io_commitROBEntries_1_ard = rob_26_ard;
        _zz_io_commitROBEntries_1_prd = rob_26_prd;
        _zz_io_commitROBEntries_1_pprd = rob_26_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_26_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_26_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_26_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_26_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_26_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_26_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_26_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_26_valid;
      end
      5'b11011 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_27_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_27_pc;
        _zz_io_commitROBEntries_1_ard = rob_27_ard;
        _zz_io_commitROBEntries_1_prd = rob_27_prd;
        _zz_io_commitROBEntries_1_pprd = rob_27_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_27_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_27_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_27_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_27_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_27_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_27_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_27_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_27_valid;
      end
      5'b11100 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_28_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_28_pc;
        _zz_io_commitROBEntries_1_ard = rob_28_ard;
        _zz_io_commitROBEntries_1_prd = rob_28_prd;
        _zz_io_commitROBEntries_1_pprd = rob_28_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_28_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_28_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_28_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_28_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_28_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_28_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_28_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_28_valid;
      end
      5'b11101 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_29_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_29_pc;
        _zz_io_commitROBEntries_1_ard = rob_29_ard;
        _zz_io_commitROBEntries_1_prd = rob_29_prd;
        _zz_io_commitROBEntries_1_pprd = rob_29_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_29_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_29_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_29_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_29_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_29_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_29_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_29_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_29_valid;
      end
      5'b11110 : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_30_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_30_pc;
        _zz_io_commitROBEntries_1_ard = rob_30_ard;
        _zz_io_commitROBEntries_1_prd = rob_30_prd;
        _zz_io_commitROBEntries_1_pprd = rob_30_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_30_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_30_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_30_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_30_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_30_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_30_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_30_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_30_valid;
      end
      default : begin
        _zz__zz_io_commitROBEntries_1_specialOp = rob_31_specialOp;
        _zz_io_commitROBEntries_1_pc_1 = rob_31_pc;
        _zz_io_commitROBEntries_1_ard = rob_31_ard;
        _zz_io_commitROBEntries_1_prd = rob_31_prd;
        _zz_io_commitROBEntries_1_pprd = rob_31_pprd;
        _zz_io_commitROBEntries_1_isComplete = rob_31_isComplete;
        _zz_io_commitROBEntries_1_branchResult_targetPC = rob_31_branchResult_targetPC;
        _zz_io_commitROBEntries_1_branchResult_branchResult = rob_31_branchResult_branchResult;
        _zz_io_commitROBEntries_1_branchResult_predictFail = rob_31_branchResult_predictFail;
        _zz_io_commitROBEntries_1_exceptionInfo_exception = rob_31_exceptionInfo_exception;
        _zz_io_commitROBEntries_1_exceptionInfo_eCode = rob_31_exceptionInfo_eCode;
        _zz_io_commitROBEntries_1_exceptionInfo_eSubCode = rob_31_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_1_valid = rob_31_valid;
      end
    endcase
  end

  always @(*) begin
    case(_zz_io_commitROBEntries_2_pc)
      5'b00000 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_0_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_0_pc;
        _zz_io_commitROBEntries_2_ard = rob_0_ard;
        _zz_io_commitROBEntries_2_prd = rob_0_prd;
        _zz_io_commitROBEntries_2_pprd = rob_0_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_0_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_0_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_0_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_0_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_0_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_0_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_0_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_0_valid;
      end
      5'b00001 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_1_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_1_pc;
        _zz_io_commitROBEntries_2_ard = rob_1_ard;
        _zz_io_commitROBEntries_2_prd = rob_1_prd;
        _zz_io_commitROBEntries_2_pprd = rob_1_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_1_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_1_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_1_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_1_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_1_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_1_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_1_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_1_valid;
      end
      5'b00010 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_2_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_2_pc;
        _zz_io_commitROBEntries_2_ard = rob_2_ard;
        _zz_io_commitROBEntries_2_prd = rob_2_prd;
        _zz_io_commitROBEntries_2_pprd = rob_2_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_2_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_2_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_2_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_2_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_2_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_2_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_2_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_2_valid;
      end
      5'b00011 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_3_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_3_pc;
        _zz_io_commitROBEntries_2_ard = rob_3_ard;
        _zz_io_commitROBEntries_2_prd = rob_3_prd;
        _zz_io_commitROBEntries_2_pprd = rob_3_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_3_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_3_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_3_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_3_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_3_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_3_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_3_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_3_valid;
      end
      5'b00100 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_4_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_4_pc;
        _zz_io_commitROBEntries_2_ard = rob_4_ard;
        _zz_io_commitROBEntries_2_prd = rob_4_prd;
        _zz_io_commitROBEntries_2_pprd = rob_4_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_4_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_4_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_4_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_4_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_4_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_4_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_4_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_4_valid;
      end
      5'b00101 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_5_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_5_pc;
        _zz_io_commitROBEntries_2_ard = rob_5_ard;
        _zz_io_commitROBEntries_2_prd = rob_5_prd;
        _zz_io_commitROBEntries_2_pprd = rob_5_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_5_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_5_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_5_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_5_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_5_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_5_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_5_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_5_valid;
      end
      5'b00110 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_6_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_6_pc;
        _zz_io_commitROBEntries_2_ard = rob_6_ard;
        _zz_io_commitROBEntries_2_prd = rob_6_prd;
        _zz_io_commitROBEntries_2_pprd = rob_6_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_6_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_6_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_6_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_6_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_6_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_6_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_6_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_6_valid;
      end
      5'b00111 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_7_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_7_pc;
        _zz_io_commitROBEntries_2_ard = rob_7_ard;
        _zz_io_commitROBEntries_2_prd = rob_7_prd;
        _zz_io_commitROBEntries_2_pprd = rob_7_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_7_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_7_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_7_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_7_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_7_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_7_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_7_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_7_valid;
      end
      5'b01000 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_8_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_8_pc;
        _zz_io_commitROBEntries_2_ard = rob_8_ard;
        _zz_io_commitROBEntries_2_prd = rob_8_prd;
        _zz_io_commitROBEntries_2_pprd = rob_8_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_8_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_8_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_8_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_8_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_8_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_8_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_8_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_8_valid;
      end
      5'b01001 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_9_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_9_pc;
        _zz_io_commitROBEntries_2_ard = rob_9_ard;
        _zz_io_commitROBEntries_2_prd = rob_9_prd;
        _zz_io_commitROBEntries_2_pprd = rob_9_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_9_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_9_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_9_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_9_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_9_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_9_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_9_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_9_valid;
      end
      5'b01010 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_10_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_10_pc;
        _zz_io_commitROBEntries_2_ard = rob_10_ard;
        _zz_io_commitROBEntries_2_prd = rob_10_prd;
        _zz_io_commitROBEntries_2_pprd = rob_10_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_10_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_10_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_10_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_10_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_10_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_10_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_10_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_10_valid;
      end
      5'b01011 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_11_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_11_pc;
        _zz_io_commitROBEntries_2_ard = rob_11_ard;
        _zz_io_commitROBEntries_2_prd = rob_11_prd;
        _zz_io_commitROBEntries_2_pprd = rob_11_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_11_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_11_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_11_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_11_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_11_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_11_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_11_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_11_valid;
      end
      5'b01100 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_12_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_12_pc;
        _zz_io_commitROBEntries_2_ard = rob_12_ard;
        _zz_io_commitROBEntries_2_prd = rob_12_prd;
        _zz_io_commitROBEntries_2_pprd = rob_12_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_12_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_12_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_12_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_12_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_12_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_12_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_12_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_12_valid;
      end
      5'b01101 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_13_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_13_pc;
        _zz_io_commitROBEntries_2_ard = rob_13_ard;
        _zz_io_commitROBEntries_2_prd = rob_13_prd;
        _zz_io_commitROBEntries_2_pprd = rob_13_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_13_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_13_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_13_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_13_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_13_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_13_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_13_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_13_valid;
      end
      5'b01110 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_14_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_14_pc;
        _zz_io_commitROBEntries_2_ard = rob_14_ard;
        _zz_io_commitROBEntries_2_prd = rob_14_prd;
        _zz_io_commitROBEntries_2_pprd = rob_14_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_14_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_14_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_14_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_14_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_14_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_14_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_14_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_14_valid;
      end
      5'b01111 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_15_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_15_pc;
        _zz_io_commitROBEntries_2_ard = rob_15_ard;
        _zz_io_commitROBEntries_2_prd = rob_15_prd;
        _zz_io_commitROBEntries_2_pprd = rob_15_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_15_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_15_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_15_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_15_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_15_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_15_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_15_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_15_valid;
      end
      5'b10000 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_16_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_16_pc;
        _zz_io_commitROBEntries_2_ard = rob_16_ard;
        _zz_io_commitROBEntries_2_prd = rob_16_prd;
        _zz_io_commitROBEntries_2_pprd = rob_16_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_16_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_16_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_16_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_16_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_16_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_16_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_16_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_16_valid;
      end
      5'b10001 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_17_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_17_pc;
        _zz_io_commitROBEntries_2_ard = rob_17_ard;
        _zz_io_commitROBEntries_2_prd = rob_17_prd;
        _zz_io_commitROBEntries_2_pprd = rob_17_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_17_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_17_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_17_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_17_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_17_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_17_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_17_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_17_valid;
      end
      5'b10010 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_18_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_18_pc;
        _zz_io_commitROBEntries_2_ard = rob_18_ard;
        _zz_io_commitROBEntries_2_prd = rob_18_prd;
        _zz_io_commitROBEntries_2_pprd = rob_18_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_18_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_18_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_18_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_18_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_18_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_18_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_18_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_18_valid;
      end
      5'b10011 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_19_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_19_pc;
        _zz_io_commitROBEntries_2_ard = rob_19_ard;
        _zz_io_commitROBEntries_2_prd = rob_19_prd;
        _zz_io_commitROBEntries_2_pprd = rob_19_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_19_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_19_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_19_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_19_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_19_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_19_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_19_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_19_valid;
      end
      5'b10100 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_20_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_20_pc;
        _zz_io_commitROBEntries_2_ard = rob_20_ard;
        _zz_io_commitROBEntries_2_prd = rob_20_prd;
        _zz_io_commitROBEntries_2_pprd = rob_20_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_20_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_20_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_20_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_20_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_20_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_20_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_20_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_20_valid;
      end
      5'b10101 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_21_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_21_pc;
        _zz_io_commitROBEntries_2_ard = rob_21_ard;
        _zz_io_commitROBEntries_2_prd = rob_21_prd;
        _zz_io_commitROBEntries_2_pprd = rob_21_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_21_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_21_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_21_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_21_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_21_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_21_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_21_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_21_valid;
      end
      5'b10110 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_22_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_22_pc;
        _zz_io_commitROBEntries_2_ard = rob_22_ard;
        _zz_io_commitROBEntries_2_prd = rob_22_prd;
        _zz_io_commitROBEntries_2_pprd = rob_22_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_22_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_22_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_22_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_22_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_22_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_22_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_22_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_22_valid;
      end
      5'b10111 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_23_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_23_pc;
        _zz_io_commitROBEntries_2_ard = rob_23_ard;
        _zz_io_commitROBEntries_2_prd = rob_23_prd;
        _zz_io_commitROBEntries_2_pprd = rob_23_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_23_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_23_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_23_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_23_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_23_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_23_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_23_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_23_valid;
      end
      5'b11000 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_24_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_24_pc;
        _zz_io_commitROBEntries_2_ard = rob_24_ard;
        _zz_io_commitROBEntries_2_prd = rob_24_prd;
        _zz_io_commitROBEntries_2_pprd = rob_24_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_24_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_24_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_24_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_24_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_24_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_24_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_24_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_24_valid;
      end
      5'b11001 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_25_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_25_pc;
        _zz_io_commitROBEntries_2_ard = rob_25_ard;
        _zz_io_commitROBEntries_2_prd = rob_25_prd;
        _zz_io_commitROBEntries_2_pprd = rob_25_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_25_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_25_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_25_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_25_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_25_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_25_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_25_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_25_valid;
      end
      5'b11010 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_26_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_26_pc;
        _zz_io_commitROBEntries_2_ard = rob_26_ard;
        _zz_io_commitROBEntries_2_prd = rob_26_prd;
        _zz_io_commitROBEntries_2_pprd = rob_26_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_26_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_26_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_26_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_26_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_26_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_26_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_26_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_26_valid;
      end
      5'b11011 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_27_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_27_pc;
        _zz_io_commitROBEntries_2_ard = rob_27_ard;
        _zz_io_commitROBEntries_2_prd = rob_27_prd;
        _zz_io_commitROBEntries_2_pprd = rob_27_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_27_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_27_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_27_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_27_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_27_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_27_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_27_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_27_valid;
      end
      5'b11100 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_28_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_28_pc;
        _zz_io_commitROBEntries_2_ard = rob_28_ard;
        _zz_io_commitROBEntries_2_prd = rob_28_prd;
        _zz_io_commitROBEntries_2_pprd = rob_28_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_28_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_28_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_28_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_28_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_28_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_28_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_28_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_28_valid;
      end
      5'b11101 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_29_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_29_pc;
        _zz_io_commitROBEntries_2_ard = rob_29_ard;
        _zz_io_commitROBEntries_2_prd = rob_29_prd;
        _zz_io_commitROBEntries_2_pprd = rob_29_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_29_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_29_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_29_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_29_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_29_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_29_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_29_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_29_valid;
      end
      5'b11110 : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_30_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_30_pc;
        _zz_io_commitROBEntries_2_ard = rob_30_ard;
        _zz_io_commitROBEntries_2_prd = rob_30_prd;
        _zz_io_commitROBEntries_2_pprd = rob_30_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_30_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_30_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_30_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_30_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_30_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_30_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_30_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_30_valid;
      end
      default : begin
        _zz__zz_io_commitROBEntries_2_specialOp = rob_31_specialOp;
        _zz_io_commitROBEntries_2_pc_1 = rob_31_pc;
        _zz_io_commitROBEntries_2_ard = rob_31_ard;
        _zz_io_commitROBEntries_2_prd = rob_31_prd;
        _zz_io_commitROBEntries_2_pprd = rob_31_pprd;
        _zz_io_commitROBEntries_2_isComplete = rob_31_isComplete;
        _zz_io_commitROBEntries_2_branchResult_targetPC = rob_31_branchResult_targetPC;
        _zz_io_commitROBEntries_2_branchResult_branchResult = rob_31_branchResult_branchResult;
        _zz_io_commitROBEntries_2_branchResult_predictFail = rob_31_branchResult_predictFail;
        _zz_io_commitROBEntries_2_exceptionInfo_exception = rob_31_exceptionInfo_exception;
        _zz_io_commitROBEntries_2_exceptionInfo_eCode = rob_31_exceptionInfo_eCode;
        _zz_io_commitROBEntries_2_exceptionInfo_eSubCode = rob_31_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_2_valid = rob_31_valid;
      end
    endcase
  end

  always @(*) begin
    case(_zz_io_commitROBEntries_3_pc)
      5'b00000 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_0_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_0_pc;
        _zz_io_commitROBEntries_3_ard = rob_0_ard;
        _zz_io_commitROBEntries_3_prd = rob_0_prd;
        _zz_io_commitROBEntries_3_pprd = rob_0_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_0_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_0_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_0_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_0_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_0_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_0_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_0_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_0_valid;
      end
      5'b00001 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_1_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_1_pc;
        _zz_io_commitROBEntries_3_ard = rob_1_ard;
        _zz_io_commitROBEntries_3_prd = rob_1_prd;
        _zz_io_commitROBEntries_3_pprd = rob_1_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_1_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_1_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_1_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_1_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_1_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_1_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_1_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_1_valid;
      end
      5'b00010 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_2_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_2_pc;
        _zz_io_commitROBEntries_3_ard = rob_2_ard;
        _zz_io_commitROBEntries_3_prd = rob_2_prd;
        _zz_io_commitROBEntries_3_pprd = rob_2_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_2_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_2_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_2_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_2_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_2_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_2_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_2_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_2_valid;
      end
      5'b00011 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_3_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_3_pc;
        _zz_io_commitROBEntries_3_ard = rob_3_ard;
        _zz_io_commitROBEntries_3_prd = rob_3_prd;
        _zz_io_commitROBEntries_3_pprd = rob_3_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_3_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_3_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_3_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_3_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_3_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_3_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_3_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_3_valid;
      end
      5'b00100 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_4_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_4_pc;
        _zz_io_commitROBEntries_3_ard = rob_4_ard;
        _zz_io_commitROBEntries_3_prd = rob_4_prd;
        _zz_io_commitROBEntries_3_pprd = rob_4_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_4_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_4_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_4_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_4_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_4_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_4_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_4_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_4_valid;
      end
      5'b00101 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_5_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_5_pc;
        _zz_io_commitROBEntries_3_ard = rob_5_ard;
        _zz_io_commitROBEntries_3_prd = rob_5_prd;
        _zz_io_commitROBEntries_3_pprd = rob_5_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_5_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_5_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_5_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_5_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_5_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_5_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_5_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_5_valid;
      end
      5'b00110 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_6_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_6_pc;
        _zz_io_commitROBEntries_3_ard = rob_6_ard;
        _zz_io_commitROBEntries_3_prd = rob_6_prd;
        _zz_io_commitROBEntries_3_pprd = rob_6_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_6_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_6_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_6_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_6_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_6_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_6_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_6_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_6_valid;
      end
      5'b00111 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_7_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_7_pc;
        _zz_io_commitROBEntries_3_ard = rob_7_ard;
        _zz_io_commitROBEntries_3_prd = rob_7_prd;
        _zz_io_commitROBEntries_3_pprd = rob_7_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_7_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_7_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_7_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_7_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_7_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_7_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_7_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_7_valid;
      end
      5'b01000 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_8_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_8_pc;
        _zz_io_commitROBEntries_3_ard = rob_8_ard;
        _zz_io_commitROBEntries_3_prd = rob_8_prd;
        _zz_io_commitROBEntries_3_pprd = rob_8_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_8_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_8_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_8_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_8_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_8_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_8_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_8_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_8_valid;
      end
      5'b01001 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_9_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_9_pc;
        _zz_io_commitROBEntries_3_ard = rob_9_ard;
        _zz_io_commitROBEntries_3_prd = rob_9_prd;
        _zz_io_commitROBEntries_3_pprd = rob_9_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_9_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_9_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_9_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_9_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_9_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_9_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_9_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_9_valid;
      end
      5'b01010 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_10_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_10_pc;
        _zz_io_commitROBEntries_3_ard = rob_10_ard;
        _zz_io_commitROBEntries_3_prd = rob_10_prd;
        _zz_io_commitROBEntries_3_pprd = rob_10_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_10_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_10_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_10_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_10_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_10_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_10_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_10_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_10_valid;
      end
      5'b01011 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_11_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_11_pc;
        _zz_io_commitROBEntries_3_ard = rob_11_ard;
        _zz_io_commitROBEntries_3_prd = rob_11_prd;
        _zz_io_commitROBEntries_3_pprd = rob_11_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_11_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_11_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_11_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_11_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_11_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_11_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_11_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_11_valid;
      end
      5'b01100 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_12_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_12_pc;
        _zz_io_commitROBEntries_3_ard = rob_12_ard;
        _zz_io_commitROBEntries_3_prd = rob_12_prd;
        _zz_io_commitROBEntries_3_pprd = rob_12_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_12_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_12_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_12_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_12_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_12_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_12_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_12_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_12_valid;
      end
      5'b01101 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_13_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_13_pc;
        _zz_io_commitROBEntries_3_ard = rob_13_ard;
        _zz_io_commitROBEntries_3_prd = rob_13_prd;
        _zz_io_commitROBEntries_3_pprd = rob_13_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_13_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_13_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_13_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_13_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_13_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_13_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_13_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_13_valid;
      end
      5'b01110 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_14_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_14_pc;
        _zz_io_commitROBEntries_3_ard = rob_14_ard;
        _zz_io_commitROBEntries_3_prd = rob_14_prd;
        _zz_io_commitROBEntries_3_pprd = rob_14_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_14_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_14_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_14_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_14_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_14_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_14_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_14_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_14_valid;
      end
      5'b01111 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_15_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_15_pc;
        _zz_io_commitROBEntries_3_ard = rob_15_ard;
        _zz_io_commitROBEntries_3_prd = rob_15_prd;
        _zz_io_commitROBEntries_3_pprd = rob_15_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_15_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_15_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_15_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_15_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_15_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_15_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_15_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_15_valid;
      end
      5'b10000 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_16_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_16_pc;
        _zz_io_commitROBEntries_3_ard = rob_16_ard;
        _zz_io_commitROBEntries_3_prd = rob_16_prd;
        _zz_io_commitROBEntries_3_pprd = rob_16_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_16_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_16_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_16_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_16_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_16_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_16_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_16_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_16_valid;
      end
      5'b10001 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_17_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_17_pc;
        _zz_io_commitROBEntries_3_ard = rob_17_ard;
        _zz_io_commitROBEntries_3_prd = rob_17_prd;
        _zz_io_commitROBEntries_3_pprd = rob_17_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_17_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_17_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_17_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_17_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_17_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_17_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_17_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_17_valid;
      end
      5'b10010 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_18_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_18_pc;
        _zz_io_commitROBEntries_3_ard = rob_18_ard;
        _zz_io_commitROBEntries_3_prd = rob_18_prd;
        _zz_io_commitROBEntries_3_pprd = rob_18_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_18_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_18_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_18_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_18_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_18_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_18_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_18_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_18_valid;
      end
      5'b10011 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_19_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_19_pc;
        _zz_io_commitROBEntries_3_ard = rob_19_ard;
        _zz_io_commitROBEntries_3_prd = rob_19_prd;
        _zz_io_commitROBEntries_3_pprd = rob_19_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_19_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_19_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_19_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_19_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_19_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_19_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_19_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_19_valid;
      end
      5'b10100 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_20_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_20_pc;
        _zz_io_commitROBEntries_3_ard = rob_20_ard;
        _zz_io_commitROBEntries_3_prd = rob_20_prd;
        _zz_io_commitROBEntries_3_pprd = rob_20_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_20_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_20_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_20_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_20_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_20_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_20_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_20_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_20_valid;
      end
      5'b10101 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_21_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_21_pc;
        _zz_io_commitROBEntries_3_ard = rob_21_ard;
        _zz_io_commitROBEntries_3_prd = rob_21_prd;
        _zz_io_commitROBEntries_3_pprd = rob_21_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_21_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_21_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_21_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_21_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_21_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_21_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_21_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_21_valid;
      end
      5'b10110 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_22_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_22_pc;
        _zz_io_commitROBEntries_3_ard = rob_22_ard;
        _zz_io_commitROBEntries_3_prd = rob_22_prd;
        _zz_io_commitROBEntries_3_pprd = rob_22_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_22_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_22_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_22_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_22_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_22_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_22_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_22_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_22_valid;
      end
      5'b10111 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_23_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_23_pc;
        _zz_io_commitROBEntries_3_ard = rob_23_ard;
        _zz_io_commitROBEntries_3_prd = rob_23_prd;
        _zz_io_commitROBEntries_3_pprd = rob_23_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_23_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_23_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_23_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_23_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_23_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_23_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_23_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_23_valid;
      end
      5'b11000 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_24_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_24_pc;
        _zz_io_commitROBEntries_3_ard = rob_24_ard;
        _zz_io_commitROBEntries_3_prd = rob_24_prd;
        _zz_io_commitROBEntries_3_pprd = rob_24_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_24_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_24_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_24_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_24_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_24_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_24_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_24_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_24_valid;
      end
      5'b11001 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_25_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_25_pc;
        _zz_io_commitROBEntries_3_ard = rob_25_ard;
        _zz_io_commitROBEntries_3_prd = rob_25_prd;
        _zz_io_commitROBEntries_3_pprd = rob_25_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_25_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_25_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_25_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_25_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_25_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_25_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_25_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_25_valid;
      end
      5'b11010 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_26_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_26_pc;
        _zz_io_commitROBEntries_3_ard = rob_26_ard;
        _zz_io_commitROBEntries_3_prd = rob_26_prd;
        _zz_io_commitROBEntries_3_pprd = rob_26_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_26_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_26_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_26_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_26_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_26_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_26_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_26_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_26_valid;
      end
      5'b11011 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_27_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_27_pc;
        _zz_io_commitROBEntries_3_ard = rob_27_ard;
        _zz_io_commitROBEntries_3_prd = rob_27_prd;
        _zz_io_commitROBEntries_3_pprd = rob_27_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_27_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_27_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_27_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_27_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_27_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_27_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_27_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_27_valid;
      end
      5'b11100 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_28_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_28_pc;
        _zz_io_commitROBEntries_3_ard = rob_28_ard;
        _zz_io_commitROBEntries_3_prd = rob_28_prd;
        _zz_io_commitROBEntries_3_pprd = rob_28_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_28_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_28_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_28_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_28_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_28_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_28_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_28_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_28_valid;
      end
      5'b11101 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_29_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_29_pc;
        _zz_io_commitROBEntries_3_ard = rob_29_ard;
        _zz_io_commitROBEntries_3_prd = rob_29_prd;
        _zz_io_commitROBEntries_3_pprd = rob_29_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_29_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_29_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_29_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_29_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_29_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_29_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_29_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_29_valid;
      end
      5'b11110 : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_30_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_30_pc;
        _zz_io_commitROBEntries_3_ard = rob_30_ard;
        _zz_io_commitROBEntries_3_prd = rob_30_prd;
        _zz_io_commitROBEntries_3_pprd = rob_30_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_30_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_30_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_30_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_30_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_30_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_30_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_30_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_30_valid;
      end
      default : begin
        _zz__zz_io_commitROBEntries_3_specialOp = rob_31_specialOp;
        _zz_io_commitROBEntries_3_pc_1 = rob_31_pc;
        _zz_io_commitROBEntries_3_ard = rob_31_ard;
        _zz_io_commitROBEntries_3_prd = rob_31_prd;
        _zz_io_commitROBEntries_3_pprd = rob_31_pprd;
        _zz_io_commitROBEntries_3_isComplete = rob_31_isComplete;
        _zz_io_commitROBEntries_3_branchResult_targetPC = rob_31_branchResult_targetPC;
        _zz_io_commitROBEntries_3_branchResult_branchResult = rob_31_branchResult_branchResult;
        _zz_io_commitROBEntries_3_branchResult_predictFail = rob_31_branchResult_predictFail;
        _zz_io_commitROBEntries_3_exceptionInfo_exception = rob_31_exceptionInfo_exception;
        _zz_io_commitROBEntries_3_exceptionInfo_eCode = rob_31_exceptionInfo_eCode;
        _zz_io_commitROBEntries_3_exceptionInfo_eSubCode = rob_31_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_3_valid = rob_31_valid;
      end
    endcase
  end

  always @(*) begin
    case(_zz_io_commitROBEntries_4_pc)
      5'b00000 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_0_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_0_pc;
        _zz_io_commitROBEntries_4_ard = rob_0_ard;
        _zz_io_commitROBEntries_4_prd = rob_0_prd;
        _zz_io_commitROBEntries_4_pprd = rob_0_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_0_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_0_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_0_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_0_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_0_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_0_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_0_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_0_valid;
      end
      5'b00001 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_1_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_1_pc;
        _zz_io_commitROBEntries_4_ard = rob_1_ard;
        _zz_io_commitROBEntries_4_prd = rob_1_prd;
        _zz_io_commitROBEntries_4_pprd = rob_1_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_1_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_1_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_1_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_1_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_1_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_1_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_1_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_1_valid;
      end
      5'b00010 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_2_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_2_pc;
        _zz_io_commitROBEntries_4_ard = rob_2_ard;
        _zz_io_commitROBEntries_4_prd = rob_2_prd;
        _zz_io_commitROBEntries_4_pprd = rob_2_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_2_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_2_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_2_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_2_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_2_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_2_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_2_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_2_valid;
      end
      5'b00011 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_3_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_3_pc;
        _zz_io_commitROBEntries_4_ard = rob_3_ard;
        _zz_io_commitROBEntries_4_prd = rob_3_prd;
        _zz_io_commitROBEntries_4_pprd = rob_3_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_3_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_3_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_3_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_3_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_3_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_3_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_3_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_3_valid;
      end
      5'b00100 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_4_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_4_pc;
        _zz_io_commitROBEntries_4_ard = rob_4_ard;
        _zz_io_commitROBEntries_4_prd = rob_4_prd;
        _zz_io_commitROBEntries_4_pprd = rob_4_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_4_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_4_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_4_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_4_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_4_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_4_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_4_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_4_valid;
      end
      5'b00101 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_5_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_5_pc;
        _zz_io_commitROBEntries_4_ard = rob_5_ard;
        _zz_io_commitROBEntries_4_prd = rob_5_prd;
        _zz_io_commitROBEntries_4_pprd = rob_5_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_5_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_5_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_5_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_5_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_5_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_5_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_5_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_5_valid;
      end
      5'b00110 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_6_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_6_pc;
        _zz_io_commitROBEntries_4_ard = rob_6_ard;
        _zz_io_commitROBEntries_4_prd = rob_6_prd;
        _zz_io_commitROBEntries_4_pprd = rob_6_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_6_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_6_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_6_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_6_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_6_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_6_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_6_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_6_valid;
      end
      5'b00111 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_7_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_7_pc;
        _zz_io_commitROBEntries_4_ard = rob_7_ard;
        _zz_io_commitROBEntries_4_prd = rob_7_prd;
        _zz_io_commitROBEntries_4_pprd = rob_7_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_7_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_7_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_7_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_7_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_7_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_7_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_7_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_7_valid;
      end
      5'b01000 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_8_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_8_pc;
        _zz_io_commitROBEntries_4_ard = rob_8_ard;
        _zz_io_commitROBEntries_4_prd = rob_8_prd;
        _zz_io_commitROBEntries_4_pprd = rob_8_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_8_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_8_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_8_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_8_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_8_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_8_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_8_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_8_valid;
      end
      5'b01001 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_9_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_9_pc;
        _zz_io_commitROBEntries_4_ard = rob_9_ard;
        _zz_io_commitROBEntries_4_prd = rob_9_prd;
        _zz_io_commitROBEntries_4_pprd = rob_9_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_9_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_9_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_9_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_9_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_9_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_9_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_9_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_9_valid;
      end
      5'b01010 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_10_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_10_pc;
        _zz_io_commitROBEntries_4_ard = rob_10_ard;
        _zz_io_commitROBEntries_4_prd = rob_10_prd;
        _zz_io_commitROBEntries_4_pprd = rob_10_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_10_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_10_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_10_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_10_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_10_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_10_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_10_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_10_valid;
      end
      5'b01011 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_11_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_11_pc;
        _zz_io_commitROBEntries_4_ard = rob_11_ard;
        _zz_io_commitROBEntries_4_prd = rob_11_prd;
        _zz_io_commitROBEntries_4_pprd = rob_11_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_11_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_11_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_11_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_11_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_11_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_11_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_11_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_11_valid;
      end
      5'b01100 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_12_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_12_pc;
        _zz_io_commitROBEntries_4_ard = rob_12_ard;
        _zz_io_commitROBEntries_4_prd = rob_12_prd;
        _zz_io_commitROBEntries_4_pprd = rob_12_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_12_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_12_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_12_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_12_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_12_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_12_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_12_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_12_valid;
      end
      5'b01101 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_13_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_13_pc;
        _zz_io_commitROBEntries_4_ard = rob_13_ard;
        _zz_io_commitROBEntries_4_prd = rob_13_prd;
        _zz_io_commitROBEntries_4_pprd = rob_13_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_13_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_13_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_13_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_13_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_13_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_13_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_13_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_13_valid;
      end
      5'b01110 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_14_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_14_pc;
        _zz_io_commitROBEntries_4_ard = rob_14_ard;
        _zz_io_commitROBEntries_4_prd = rob_14_prd;
        _zz_io_commitROBEntries_4_pprd = rob_14_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_14_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_14_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_14_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_14_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_14_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_14_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_14_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_14_valid;
      end
      5'b01111 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_15_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_15_pc;
        _zz_io_commitROBEntries_4_ard = rob_15_ard;
        _zz_io_commitROBEntries_4_prd = rob_15_prd;
        _zz_io_commitROBEntries_4_pprd = rob_15_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_15_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_15_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_15_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_15_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_15_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_15_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_15_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_15_valid;
      end
      5'b10000 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_16_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_16_pc;
        _zz_io_commitROBEntries_4_ard = rob_16_ard;
        _zz_io_commitROBEntries_4_prd = rob_16_prd;
        _zz_io_commitROBEntries_4_pprd = rob_16_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_16_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_16_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_16_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_16_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_16_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_16_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_16_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_16_valid;
      end
      5'b10001 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_17_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_17_pc;
        _zz_io_commitROBEntries_4_ard = rob_17_ard;
        _zz_io_commitROBEntries_4_prd = rob_17_prd;
        _zz_io_commitROBEntries_4_pprd = rob_17_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_17_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_17_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_17_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_17_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_17_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_17_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_17_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_17_valid;
      end
      5'b10010 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_18_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_18_pc;
        _zz_io_commitROBEntries_4_ard = rob_18_ard;
        _zz_io_commitROBEntries_4_prd = rob_18_prd;
        _zz_io_commitROBEntries_4_pprd = rob_18_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_18_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_18_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_18_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_18_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_18_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_18_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_18_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_18_valid;
      end
      5'b10011 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_19_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_19_pc;
        _zz_io_commitROBEntries_4_ard = rob_19_ard;
        _zz_io_commitROBEntries_4_prd = rob_19_prd;
        _zz_io_commitROBEntries_4_pprd = rob_19_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_19_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_19_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_19_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_19_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_19_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_19_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_19_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_19_valid;
      end
      5'b10100 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_20_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_20_pc;
        _zz_io_commitROBEntries_4_ard = rob_20_ard;
        _zz_io_commitROBEntries_4_prd = rob_20_prd;
        _zz_io_commitROBEntries_4_pprd = rob_20_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_20_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_20_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_20_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_20_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_20_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_20_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_20_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_20_valid;
      end
      5'b10101 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_21_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_21_pc;
        _zz_io_commitROBEntries_4_ard = rob_21_ard;
        _zz_io_commitROBEntries_4_prd = rob_21_prd;
        _zz_io_commitROBEntries_4_pprd = rob_21_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_21_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_21_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_21_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_21_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_21_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_21_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_21_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_21_valid;
      end
      5'b10110 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_22_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_22_pc;
        _zz_io_commitROBEntries_4_ard = rob_22_ard;
        _zz_io_commitROBEntries_4_prd = rob_22_prd;
        _zz_io_commitROBEntries_4_pprd = rob_22_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_22_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_22_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_22_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_22_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_22_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_22_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_22_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_22_valid;
      end
      5'b10111 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_23_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_23_pc;
        _zz_io_commitROBEntries_4_ard = rob_23_ard;
        _zz_io_commitROBEntries_4_prd = rob_23_prd;
        _zz_io_commitROBEntries_4_pprd = rob_23_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_23_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_23_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_23_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_23_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_23_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_23_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_23_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_23_valid;
      end
      5'b11000 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_24_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_24_pc;
        _zz_io_commitROBEntries_4_ard = rob_24_ard;
        _zz_io_commitROBEntries_4_prd = rob_24_prd;
        _zz_io_commitROBEntries_4_pprd = rob_24_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_24_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_24_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_24_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_24_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_24_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_24_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_24_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_24_valid;
      end
      5'b11001 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_25_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_25_pc;
        _zz_io_commitROBEntries_4_ard = rob_25_ard;
        _zz_io_commitROBEntries_4_prd = rob_25_prd;
        _zz_io_commitROBEntries_4_pprd = rob_25_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_25_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_25_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_25_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_25_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_25_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_25_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_25_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_25_valid;
      end
      5'b11010 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_26_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_26_pc;
        _zz_io_commitROBEntries_4_ard = rob_26_ard;
        _zz_io_commitROBEntries_4_prd = rob_26_prd;
        _zz_io_commitROBEntries_4_pprd = rob_26_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_26_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_26_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_26_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_26_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_26_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_26_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_26_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_26_valid;
      end
      5'b11011 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_27_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_27_pc;
        _zz_io_commitROBEntries_4_ard = rob_27_ard;
        _zz_io_commitROBEntries_4_prd = rob_27_prd;
        _zz_io_commitROBEntries_4_pprd = rob_27_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_27_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_27_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_27_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_27_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_27_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_27_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_27_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_27_valid;
      end
      5'b11100 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_28_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_28_pc;
        _zz_io_commitROBEntries_4_ard = rob_28_ard;
        _zz_io_commitROBEntries_4_prd = rob_28_prd;
        _zz_io_commitROBEntries_4_pprd = rob_28_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_28_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_28_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_28_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_28_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_28_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_28_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_28_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_28_valid;
      end
      5'b11101 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_29_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_29_pc;
        _zz_io_commitROBEntries_4_ard = rob_29_ard;
        _zz_io_commitROBEntries_4_prd = rob_29_prd;
        _zz_io_commitROBEntries_4_pprd = rob_29_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_29_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_29_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_29_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_29_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_29_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_29_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_29_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_29_valid;
      end
      5'b11110 : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_30_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_30_pc;
        _zz_io_commitROBEntries_4_ard = rob_30_ard;
        _zz_io_commitROBEntries_4_prd = rob_30_prd;
        _zz_io_commitROBEntries_4_pprd = rob_30_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_30_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_30_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_30_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_30_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_30_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_30_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_30_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_30_valid;
      end
      default : begin
        _zz__zz_io_commitROBEntries_4_specialOp = rob_31_specialOp;
        _zz_io_commitROBEntries_4_pc_1 = rob_31_pc;
        _zz_io_commitROBEntries_4_ard = rob_31_ard;
        _zz_io_commitROBEntries_4_prd = rob_31_prd;
        _zz_io_commitROBEntries_4_pprd = rob_31_pprd;
        _zz_io_commitROBEntries_4_isComplete = rob_31_isComplete;
        _zz_io_commitROBEntries_4_branchResult_targetPC = rob_31_branchResult_targetPC;
        _zz_io_commitROBEntries_4_branchResult_branchResult = rob_31_branchResult_branchResult;
        _zz_io_commitROBEntries_4_branchResult_predictFail = rob_31_branchResult_predictFail;
        _zz_io_commitROBEntries_4_exceptionInfo_exception = rob_31_exceptionInfo_exception;
        _zz_io_commitROBEntries_4_exceptionInfo_eCode = rob_31_exceptionInfo_eCode;
        _zz_io_commitROBEntries_4_exceptionInfo_eSubCode = rob_31_exceptionInfo_eSubCode;
        _zz_io_commitROBEntries_4_valid = rob_31_valid;
      end
    endcase
  end

  always @(*) begin
    case(_zz_stage_freePRFNum_2)
      2'b00 : _zz_stage_freePRFNum_1 = 2'b00;
      2'b01 : _zz_stage_freePRFNum_1 = 2'b01;
      2'b10 : _zz_stage_freePRFNum_1 = 2'b01;
      default : _zz_stage_freePRFNum_1 = 2'b10;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_dispatch_specialOp_0)
      ROBSpecialOp_nop : io_dispatch_specialOp_0_string = "nop      ";
      ROBSpecialOp_bpuUpdate : io_dispatch_specialOp_0_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : io_dispatch_specialOp_0_string = "lsuAction";
      ROBSpecialOp_ll : io_dispatch_specialOp_0_string = "ll       ";
      ROBSpecialOp_writeCSR : io_dispatch_specialOp_0_string = "writeCSR ";
      ROBSpecialOp_ertn : io_dispatch_specialOp_0_string = "ertn     ";
      ROBSpecialOp_idle : io_dispatch_specialOp_0_string = "idle     ";
      ROBSpecialOp_readCSR : io_dispatch_specialOp_0_string = "readCSR  ";
      ROBSpecialOp_readCNT : io_dispatch_specialOp_0_string = "readCNT  ";
      default : io_dispatch_specialOp_0_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_dispatch_specialOp_1)
      ROBSpecialOp_nop : io_dispatch_specialOp_1_string = "nop      ";
      ROBSpecialOp_bpuUpdate : io_dispatch_specialOp_1_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : io_dispatch_specialOp_1_string = "lsuAction";
      ROBSpecialOp_ll : io_dispatch_specialOp_1_string = "ll       ";
      ROBSpecialOp_writeCSR : io_dispatch_specialOp_1_string = "writeCSR ";
      ROBSpecialOp_ertn : io_dispatch_specialOp_1_string = "ertn     ";
      ROBSpecialOp_idle : io_dispatch_specialOp_1_string = "idle     ";
      ROBSpecialOp_readCSR : io_dispatch_specialOp_1_string = "readCSR  ";
      ROBSpecialOp_readCNT : io_dispatch_specialOp_1_string = "readCNT  ";
      default : io_dispatch_specialOp_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_commitROBEntries_0_specialOp)
      ROBSpecialOp_nop : io_commitROBEntries_0_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : io_commitROBEntries_0_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : io_commitROBEntries_0_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : io_commitROBEntries_0_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : io_commitROBEntries_0_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : io_commitROBEntries_0_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : io_commitROBEntries_0_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : io_commitROBEntries_0_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : io_commitROBEntries_0_specialOp_string = "readCNT  ";
      default : io_commitROBEntries_0_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_commitROBEntries_1_specialOp)
      ROBSpecialOp_nop : io_commitROBEntries_1_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : io_commitROBEntries_1_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : io_commitROBEntries_1_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : io_commitROBEntries_1_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : io_commitROBEntries_1_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : io_commitROBEntries_1_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : io_commitROBEntries_1_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : io_commitROBEntries_1_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : io_commitROBEntries_1_specialOp_string = "readCNT  ";
      default : io_commitROBEntries_1_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_commitROBEntries_2_specialOp)
      ROBSpecialOp_nop : io_commitROBEntries_2_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : io_commitROBEntries_2_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : io_commitROBEntries_2_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : io_commitROBEntries_2_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : io_commitROBEntries_2_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : io_commitROBEntries_2_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : io_commitROBEntries_2_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : io_commitROBEntries_2_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : io_commitROBEntries_2_specialOp_string = "readCNT  ";
      default : io_commitROBEntries_2_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_commitROBEntries_3_specialOp)
      ROBSpecialOp_nop : io_commitROBEntries_3_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : io_commitROBEntries_3_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : io_commitROBEntries_3_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : io_commitROBEntries_3_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : io_commitROBEntries_3_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : io_commitROBEntries_3_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : io_commitROBEntries_3_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : io_commitROBEntries_3_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : io_commitROBEntries_3_specialOp_string = "readCNT  ";
      default : io_commitROBEntries_3_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_commitROBEntries_4_specialOp)
      ROBSpecialOp_nop : io_commitROBEntries_4_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : io_commitROBEntries_4_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : io_commitROBEntries_4_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : io_commitROBEntries_4_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : io_commitROBEntries_4_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : io_commitROBEntries_4_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : io_commitROBEntries_4_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : io_commitROBEntries_4_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : io_commitROBEntries_4_specialOp_string = "readCNT  ";
      default : io_commitROBEntries_4_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_0_specialOp)
      ROBSpecialOp_nop : rob_0_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_0_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_0_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_0_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_0_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_0_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_0_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_0_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_0_specialOp_string = "readCNT  ";
      default : rob_0_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_1_specialOp)
      ROBSpecialOp_nop : rob_1_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_1_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_1_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_1_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_1_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_1_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_1_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_1_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_1_specialOp_string = "readCNT  ";
      default : rob_1_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_2_specialOp)
      ROBSpecialOp_nop : rob_2_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_2_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_2_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_2_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_2_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_2_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_2_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_2_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_2_specialOp_string = "readCNT  ";
      default : rob_2_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_3_specialOp)
      ROBSpecialOp_nop : rob_3_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_3_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_3_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_3_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_3_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_3_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_3_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_3_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_3_specialOp_string = "readCNT  ";
      default : rob_3_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_4_specialOp)
      ROBSpecialOp_nop : rob_4_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_4_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_4_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_4_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_4_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_4_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_4_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_4_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_4_specialOp_string = "readCNT  ";
      default : rob_4_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_5_specialOp)
      ROBSpecialOp_nop : rob_5_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_5_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_5_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_5_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_5_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_5_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_5_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_5_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_5_specialOp_string = "readCNT  ";
      default : rob_5_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_6_specialOp)
      ROBSpecialOp_nop : rob_6_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_6_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_6_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_6_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_6_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_6_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_6_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_6_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_6_specialOp_string = "readCNT  ";
      default : rob_6_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_7_specialOp)
      ROBSpecialOp_nop : rob_7_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_7_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_7_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_7_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_7_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_7_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_7_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_7_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_7_specialOp_string = "readCNT  ";
      default : rob_7_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_8_specialOp)
      ROBSpecialOp_nop : rob_8_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_8_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_8_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_8_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_8_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_8_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_8_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_8_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_8_specialOp_string = "readCNT  ";
      default : rob_8_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_9_specialOp)
      ROBSpecialOp_nop : rob_9_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_9_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_9_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_9_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_9_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_9_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_9_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_9_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_9_specialOp_string = "readCNT  ";
      default : rob_9_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_10_specialOp)
      ROBSpecialOp_nop : rob_10_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_10_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_10_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_10_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_10_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_10_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_10_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_10_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_10_specialOp_string = "readCNT  ";
      default : rob_10_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_11_specialOp)
      ROBSpecialOp_nop : rob_11_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_11_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_11_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_11_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_11_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_11_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_11_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_11_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_11_specialOp_string = "readCNT  ";
      default : rob_11_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_12_specialOp)
      ROBSpecialOp_nop : rob_12_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_12_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_12_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_12_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_12_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_12_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_12_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_12_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_12_specialOp_string = "readCNT  ";
      default : rob_12_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_13_specialOp)
      ROBSpecialOp_nop : rob_13_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_13_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_13_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_13_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_13_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_13_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_13_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_13_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_13_specialOp_string = "readCNT  ";
      default : rob_13_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_14_specialOp)
      ROBSpecialOp_nop : rob_14_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_14_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_14_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_14_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_14_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_14_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_14_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_14_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_14_specialOp_string = "readCNT  ";
      default : rob_14_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_15_specialOp)
      ROBSpecialOp_nop : rob_15_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_15_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_15_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_15_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_15_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_15_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_15_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_15_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_15_specialOp_string = "readCNT  ";
      default : rob_15_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_16_specialOp)
      ROBSpecialOp_nop : rob_16_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_16_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_16_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_16_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_16_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_16_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_16_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_16_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_16_specialOp_string = "readCNT  ";
      default : rob_16_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_17_specialOp)
      ROBSpecialOp_nop : rob_17_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_17_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_17_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_17_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_17_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_17_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_17_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_17_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_17_specialOp_string = "readCNT  ";
      default : rob_17_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_18_specialOp)
      ROBSpecialOp_nop : rob_18_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_18_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_18_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_18_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_18_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_18_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_18_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_18_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_18_specialOp_string = "readCNT  ";
      default : rob_18_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_19_specialOp)
      ROBSpecialOp_nop : rob_19_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_19_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_19_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_19_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_19_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_19_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_19_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_19_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_19_specialOp_string = "readCNT  ";
      default : rob_19_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_20_specialOp)
      ROBSpecialOp_nop : rob_20_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_20_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_20_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_20_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_20_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_20_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_20_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_20_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_20_specialOp_string = "readCNT  ";
      default : rob_20_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_21_specialOp)
      ROBSpecialOp_nop : rob_21_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_21_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_21_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_21_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_21_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_21_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_21_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_21_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_21_specialOp_string = "readCNT  ";
      default : rob_21_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_22_specialOp)
      ROBSpecialOp_nop : rob_22_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_22_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_22_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_22_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_22_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_22_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_22_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_22_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_22_specialOp_string = "readCNT  ";
      default : rob_22_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_23_specialOp)
      ROBSpecialOp_nop : rob_23_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_23_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_23_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_23_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_23_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_23_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_23_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_23_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_23_specialOp_string = "readCNT  ";
      default : rob_23_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_24_specialOp)
      ROBSpecialOp_nop : rob_24_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_24_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_24_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_24_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_24_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_24_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_24_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_24_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_24_specialOp_string = "readCNT  ";
      default : rob_24_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_25_specialOp)
      ROBSpecialOp_nop : rob_25_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_25_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_25_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_25_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_25_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_25_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_25_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_25_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_25_specialOp_string = "readCNT  ";
      default : rob_25_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_26_specialOp)
      ROBSpecialOp_nop : rob_26_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_26_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_26_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_26_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_26_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_26_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_26_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_26_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_26_specialOp_string = "readCNT  ";
      default : rob_26_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_27_specialOp)
      ROBSpecialOp_nop : rob_27_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_27_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_27_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_27_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_27_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_27_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_27_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_27_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_27_specialOp_string = "readCNT  ";
      default : rob_27_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_28_specialOp)
      ROBSpecialOp_nop : rob_28_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_28_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_28_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_28_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_28_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_28_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_28_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_28_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_28_specialOp_string = "readCNT  ";
      default : rob_28_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_29_specialOp)
      ROBSpecialOp_nop : rob_29_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_29_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_29_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_29_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_29_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_29_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_29_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_29_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_29_specialOp_string = "readCNT  ";
      default : rob_29_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_30_specialOp)
      ROBSpecialOp_nop : rob_30_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_30_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_30_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_30_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_30_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_30_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_30_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_30_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_30_specialOp_string = "readCNT  ";
      default : rob_30_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rob_31_specialOp)
      ROBSpecialOp_nop : rob_31_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : rob_31_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : rob_31_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : rob_31_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : rob_31_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : rob_31_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : rob_31_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : rob_31_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : rob_31_specialOp_string = "readCNT  ";
      default : rob_31_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_stage_updateBPU_0_isJumpInst)
      ROBSpecialOp_nop : _zz_stage_updateBPU_0_isJumpInst_string = "nop      ";
      ROBSpecialOp_bpuUpdate : _zz_stage_updateBPU_0_isJumpInst_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : _zz_stage_updateBPU_0_isJumpInst_string = "lsuAction";
      ROBSpecialOp_ll : _zz_stage_updateBPU_0_isJumpInst_string = "ll       ";
      ROBSpecialOp_writeCSR : _zz_stage_updateBPU_0_isJumpInst_string = "writeCSR ";
      ROBSpecialOp_ertn : _zz_stage_updateBPU_0_isJumpInst_string = "ertn     ";
      ROBSpecialOp_idle : _zz_stage_updateBPU_0_isJumpInst_string = "idle     ";
      ROBSpecialOp_readCSR : _zz_stage_updateBPU_0_isJumpInst_string = "readCSR  ";
      ROBSpecialOp_readCNT : _zz_stage_updateBPU_0_isJumpInst_string = "readCNT  ";
      default : _zz_stage_updateBPU_0_isJumpInst_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_stage_updateBPU_1_isJumpInst)
      ROBSpecialOp_nop : _zz_stage_updateBPU_1_isJumpInst_string = "nop      ";
      ROBSpecialOp_bpuUpdate : _zz_stage_updateBPU_1_isJumpInst_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : _zz_stage_updateBPU_1_isJumpInst_string = "lsuAction";
      ROBSpecialOp_ll : _zz_stage_updateBPU_1_isJumpInst_string = "ll       ";
      ROBSpecialOp_writeCSR : _zz_stage_updateBPU_1_isJumpInst_string = "writeCSR ";
      ROBSpecialOp_ertn : _zz_stage_updateBPU_1_isJumpInst_string = "ertn     ";
      ROBSpecialOp_idle : _zz_stage_updateBPU_1_isJumpInst_string = "idle     ";
      ROBSpecialOp_readCSR : _zz_stage_updateBPU_1_isJumpInst_string = "readCSR  ";
      ROBSpecialOp_readCNT : _zz_stage_updateBPU_1_isJumpInst_string = "readCNT  ";
      default : _zz_stage_updateBPU_1_isJumpInst_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commitROBEntries_0_specialOp)
      ROBSpecialOp_nop : _zz_io_commitROBEntries_0_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : _zz_io_commitROBEntries_0_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : _zz_io_commitROBEntries_0_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : _zz_io_commitROBEntries_0_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : _zz_io_commitROBEntries_0_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : _zz_io_commitROBEntries_0_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : _zz_io_commitROBEntries_0_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : _zz_io_commitROBEntries_0_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : _zz_io_commitROBEntries_0_specialOp_string = "readCNT  ";
      default : _zz_io_commitROBEntries_0_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commitROBEntries_1_specialOp)
      ROBSpecialOp_nop : _zz_io_commitROBEntries_1_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : _zz_io_commitROBEntries_1_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : _zz_io_commitROBEntries_1_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : _zz_io_commitROBEntries_1_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : _zz_io_commitROBEntries_1_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : _zz_io_commitROBEntries_1_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : _zz_io_commitROBEntries_1_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : _zz_io_commitROBEntries_1_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : _zz_io_commitROBEntries_1_specialOp_string = "readCNT  ";
      default : _zz_io_commitROBEntries_1_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commitROBEntries_2_specialOp)
      ROBSpecialOp_nop : _zz_io_commitROBEntries_2_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : _zz_io_commitROBEntries_2_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : _zz_io_commitROBEntries_2_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : _zz_io_commitROBEntries_2_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : _zz_io_commitROBEntries_2_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : _zz_io_commitROBEntries_2_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : _zz_io_commitROBEntries_2_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : _zz_io_commitROBEntries_2_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : _zz_io_commitROBEntries_2_specialOp_string = "readCNT  ";
      default : _zz_io_commitROBEntries_2_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commitROBEntries_3_specialOp)
      ROBSpecialOp_nop : _zz_io_commitROBEntries_3_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : _zz_io_commitROBEntries_3_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : _zz_io_commitROBEntries_3_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : _zz_io_commitROBEntries_3_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : _zz_io_commitROBEntries_3_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : _zz_io_commitROBEntries_3_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : _zz_io_commitROBEntries_3_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : _zz_io_commitROBEntries_3_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : _zz_io_commitROBEntries_3_specialOp_string = "readCNT  ";
      default : _zz_io_commitROBEntries_3_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_commitROBEntries_4_specialOp)
      ROBSpecialOp_nop : _zz_io_commitROBEntries_4_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : _zz_io_commitROBEntries_4_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : _zz_io_commitROBEntries_4_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : _zz_io_commitROBEntries_4_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : _zz_io_commitROBEntries_4_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : _zz_io_commitROBEntries_4_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : _zz_io_commitROBEntries_4_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : _zz_io_commitROBEntries_4_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : _zz_io_commitROBEntries_4_specialOp_string = "readCNT  ";
      default : _zz_io_commitROBEntries_4_specialOp_string = "?????????";
    endcase
  end
  `endif

  assign _zz_retirePC_0 = _zz__zz_retirePC_0;
  assign _zz_noPPRDMask = _zz__zz_noPPRDMask;
  assign _zz_stage_updateBPU_0_isJumpInst = _zz__zz_stage_updateBPU_0_isJumpInst;
  assign _zz_retireMask = _zz__zz_retireMask;
  assign _zz_stage_updateBPU_0_taken = _zz__zz_stage_updateBPU_0_taken;
  assign _zz_stage_updateBPU_0_predictFail = _zz__zz_stage_updateBPU_0_predictFail;
  assign _zz_retireMask_1 = _zz__zz_retireMask_1;
  assign _zz_normalExceptionMask = _zz__zz_normalExceptionMask;
  assign _zz_normalExceptionMask_1 = _zz__zz_normalExceptionMask_1;
  assign _zz_retireMask_2 = _zz__zz_retireMask_2;
  assign idleEn = ((_zz_retireMask_2 && (_zz_stage_updateBPU_0_isJumpInst == ROBSpecialOp_idle)) && io_interrupt);
  assign dispatchNum = _zz_dispatchNum;
  assign retireNum = _zz_retireNum;
  always @(*) begin
    stage_availROBMask[0] = (! _zz_stage_availROBMask);
    stage_availROBMask[1] = (! _zz_stage_availROBMask_3);
  end

  assign io_dispatch_robIdx_0 = tail_0;
  assign io_dispatch_robIdx_1 = tail_1;
  always @(*) begin
    retireMask[0] = ((_zz_retireMask_2 && _zz_retireMask) && (! _zz_retireMask_1));
    retireMask[1] = ((((_zz_retireMask_5 && _zz_retireMask_3) && (! _zz_retireMask_4)) && (&retireMask[0 : 0])) && (! inhibitNextRetireMask[0]));
  end

  always @(*) begin
    flushMask[0] = ((_zz_retireMask_2 && _zz_retireMask) && (_zz_retireMask_1 || inhibitNextRetireMask[0]));
    flushMask[1] = ((((_zz_retireMask_5 && _zz_retireMask_3) && (_zz_retireMask_4 || inhibitNextRetireMask[1])) && (&retireMask[0 : 0])) && (! inhibitNextRetireMask[0]));
  end

  assign _zz_retirePC_1 = _zz__zz_retirePC_1;
  assign _zz_stage_updateBPU_1_isJumpInst = _zz__zz_stage_updateBPU_1_isJumpInst;
  assign _zz_retireMask_3 = _zz__zz_retireMask_3;
  assign _zz_stage_updateBPU_1_taken = _zz__zz_stage_updateBPU_1_taken;
  assign _zz_stage_updateBPU_1_predictFail = _zz__zz_stage_updateBPU_1_predictFail;
  assign _zz_retireMask_4 = _zz__zz_retireMask_4;
  assign _zz_normalExceptionMask_2 = _zz__zz_normalExceptionMask_2;
  assign _zz_normalExceptionMask_3 = _zz__zz_normalExceptionMask_3;
  assign _zz_retireMask_5 = _zz__zz_retireMask_5;
  assign flush = ((|flushMask) || idleEn);
  always @(*) begin
    _zz_rob_0_valid[0] = ((tail_0 == 5'h00) && io_dispatch_allowMask[0]);
    _zz_rob_0_valid[1] = ((tail_1 == 5'h00) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_0_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h00));
    _zz_rob_0_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h00));
    _zz_rob_0_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h00));
    _zz_rob_0_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h00));
    _zz_rob_0_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h00));
  end

  always @(*) begin
    _zz_rob_0_isComplete_1[0] = ((head_0 == 5'h00) && retireMask[0]);
    _zz_rob_0_isComplete_1[1] = ((head_1 == 5'h00) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_1_valid[0] = ((tail_0 == 5'h01) && io_dispatch_allowMask[0]);
    _zz_rob_1_valid[1] = ((tail_1 == 5'h01) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_1_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h01));
    _zz_rob_1_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h01));
    _zz_rob_1_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h01));
    _zz_rob_1_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h01));
    _zz_rob_1_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h01));
  end

  always @(*) begin
    _zz_rob_1_isComplete_1[0] = ((head_0 == 5'h01) && retireMask[0]);
    _zz_rob_1_isComplete_1[1] = ((head_1 == 5'h01) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_2_valid[0] = ((tail_0 == 5'h02) && io_dispatch_allowMask[0]);
    _zz_rob_2_valid[1] = ((tail_1 == 5'h02) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_2_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h02));
    _zz_rob_2_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h02));
    _zz_rob_2_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h02));
    _zz_rob_2_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h02));
    _zz_rob_2_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h02));
  end

  always @(*) begin
    _zz_rob_2_isComplete_1[0] = ((head_0 == 5'h02) && retireMask[0]);
    _zz_rob_2_isComplete_1[1] = ((head_1 == 5'h02) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_3_valid[0] = ((tail_0 == 5'h03) && io_dispatch_allowMask[0]);
    _zz_rob_3_valid[1] = ((tail_1 == 5'h03) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_3_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h03));
    _zz_rob_3_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h03));
    _zz_rob_3_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h03));
    _zz_rob_3_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h03));
    _zz_rob_3_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h03));
  end

  always @(*) begin
    _zz_rob_3_isComplete_1[0] = ((head_0 == 5'h03) && retireMask[0]);
    _zz_rob_3_isComplete_1[1] = ((head_1 == 5'h03) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_4_valid[0] = ((tail_0 == 5'h04) && io_dispatch_allowMask[0]);
    _zz_rob_4_valid[1] = ((tail_1 == 5'h04) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_4_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h04));
    _zz_rob_4_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h04));
    _zz_rob_4_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h04));
    _zz_rob_4_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h04));
    _zz_rob_4_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h04));
  end

  always @(*) begin
    _zz_rob_4_isComplete_1[0] = ((head_0 == 5'h04) && retireMask[0]);
    _zz_rob_4_isComplete_1[1] = ((head_1 == 5'h04) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_5_valid[0] = ((tail_0 == 5'h05) && io_dispatch_allowMask[0]);
    _zz_rob_5_valid[1] = ((tail_1 == 5'h05) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_5_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h05));
    _zz_rob_5_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h05));
    _zz_rob_5_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h05));
    _zz_rob_5_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h05));
    _zz_rob_5_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h05));
  end

  always @(*) begin
    _zz_rob_5_isComplete_1[0] = ((head_0 == 5'h05) && retireMask[0]);
    _zz_rob_5_isComplete_1[1] = ((head_1 == 5'h05) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_6_valid[0] = ((tail_0 == 5'h06) && io_dispatch_allowMask[0]);
    _zz_rob_6_valid[1] = ((tail_1 == 5'h06) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_6_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h06));
    _zz_rob_6_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h06));
    _zz_rob_6_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h06));
    _zz_rob_6_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h06));
    _zz_rob_6_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h06));
  end

  always @(*) begin
    _zz_rob_6_isComplete_1[0] = ((head_0 == 5'h06) && retireMask[0]);
    _zz_rob_6_isComplete_1[1] = ((head_1 == 5'h06) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_7_valid[0] = ((tail_0 == 5'h07) && io_dispatch_allowMask[0]);
    _zz_rob_7_valid[1] = ((tail_1 == 5'h07) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_7_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h07));
    _zz_rob_7_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h07));
    _zz_rob_7_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h07));
    _zz_rob_7_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h07));
    _zz_rob_7_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h07));
  end

  always @(*) begin
    _zz_rob_7_isComplete_1[0] = ((head_0 == 5'h07) && retireMask[0]);
    _zz_rob_7_isComplete_1[1] = ((head_1 == 5'h07) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_8_valid[0] = ((tail_0 == 5'h08) && io_dispatch_allowMask[0]);
    _zz_rob_8_valid[1] = ((tail_1 == 5'h08) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_8_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h08));
    _zz_rob_8_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h08));
    _zz_rob_8_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h08));
    _zz_rob_8_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h08));
    _zz_rob_8_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h08));
  end

  always @(*) begin
    _zz_rob_8_isComplete_1[0] = ((head_0 == 5'h08) && retireMask[0]);
    _zz_rob_8_isComplete_1[1] = ((head_1 == 5'h08) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_9_valid[0] = ((tail_0 == 5'h09) && io_dispatch_allowMask[0]);
    _zz_rob_9_valid[1] = ((tail_1 == 5'h09) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_9_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h09));
    _zz_rob_9_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h09));
    _zz_rob_9_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h09));
    _zz_rob_9_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h09));
    _zz_rob_9_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h09));
  end

  always @(*) begin
    _zz_rob_9_isComplete_1[0] = ((head_0 == 5'h09) && retireMask[0]);
    _zz_rob_9_isComplete_1[1] = ((head_1 == 5'h09) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_10_valid[0] = ((tail_0 == 5'h0a) && io_dispatch_allowMask[0]);
    _zz_rob_10_valid[1] = ((tail_1 == 5'h0a) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_10_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h0a));
    _zz_rob_10_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h0a));
    _zz_rob_10_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h0a));
    _zz_rob_10_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h0a));
    _zz_rob_10_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h0a));
  end

  always @(*) begin
    _zz_rob_10_isComplete_1[0] = ((head_0 == 5'h0a) && retireMask[0]);
    _zz_rob_10_isComplete_1[1] = ((head_1 == 5'h0a) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_11_valid[0] = ((tail_0 == 5'h0b) && io_dispatch_allowMask[0]);
    _zz_rob_11_valid[1] = ((tail_1 == 5'h0b) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_11_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h0b));
    _zz_rob_11_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h0b));
    _zz_rob_11_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h0b));
    _zz_rob_11_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h0b));
    _zz_rob_11_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h0b));
  end

  always @(*) begin
    _zz_rob_11_isComplete_1[0] = ((head_0 == 5'h0b) && retireMask[0]);
    _zz_rob_11_isComplete_1[1] = ((head_1 == 5'h0b) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_12_valid[0] = ((tail_0 == 5'h0c) && io_dispatch_allowMask[0]);
    _zz_rob_12_valid[1] = ((tail_1 == 5'h0c) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_12_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h0c));
    _zz_rob_12_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h0c));
    _zz_rob_12_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h0c));
    _zz_rob_12_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h0c));
    _zz_rob_12_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h0c));
  end

  always @(*) begin
    _zz_rob_12_isComplete_1[0] = ((head_0 == 5'h0c) && retireMask[0]);
    _zz_rob_12_isComplete_1[1] = ((head_1 == 5'h0c) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_13_valid[0] = ((tail_0 == 5'h0d) && io_dispatch_allowMask[0]);
    _zz_rob_13_valid[1] = ((tail_1 == 5'h0d) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_13_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h0d));
    _zz_rob_13_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h0d));
    _zz_rob_13_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h0d));
    _zz_rob_13_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h0d));
    _zz_rob_13_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h0d));
  end

  always @(*) begin
    _zz_rob_13_isComplete_1[0] = ((head_0 == 5'h0d) && retireMask[0]);
    _zz_rob_13_isComplete_1[1] = ((head_1 == 5'h0d) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_14_valid[0] = ((tail_0 == 5'h0e) && io_dispatch_allowMask[0]);
    _zz_rob_14_valid[1] = ((tail_1 == 5'h0e) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_14_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h0e));
    _zz_rob_14_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h0e));
    _zz_rob_14_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h0e));
    _zz_rob_14_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h0e));
    _zz_rob_14_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h0e));
  end

  always @(*) begin
    _zz_rob_14_isComplete_1[0] = ((head_0 == 5'h0e) && retireMask[0]);
    _zz_rob_14_isComplete_1[1] = ((head_1 == 5'h0e) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_15_valid[0] = ((tail_0 == 5'h0f) && io_dispatch_allowMask[0]);
    _zz_rob_15_valid[1] = ((tail_1 == 5'h0f) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_15_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h0f));
    _zz_rob_15_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h0f));
    _zz_rob_15_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h0f));
    _zz_rob_15_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h0f));
    _zz_rob_15_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h0f));
  end

  always @(*) begin
    _zz_rob_15_isComplete_1[0] = ((head_0 == 5'h0f) && retireMask[0]);
    _zz_rob_15_isComplete_1[1] = ((head_1 == 5'h0f) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_16_valid[0] = ((tail_0 == 5'h10) && io_dispatch_allowMask[0]);
    _zz_rob_16_valid[1] = ((tail_1 == 5'h10) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_16_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h10));
    _zz_rob_16_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h10));
    _zz_rob_16_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h10));
    _zz_rob_16_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h10));
    _zz_rob_16_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h10));
  end

  always @(*) begin
    _zz_rob_16_isComplete_1[0] = ((head_0 == 5'h10) && retireMask[0]);
    _zz_rob_16_isComplete_1[1] = ((head_1 == 5'h10) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_17_valid[0] = ((tail_0 == 5'h11) && io_dispatch_allowMask[0]);
    _zz_rob_17_valid[1] = ((tail_1 == 5'h11) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_17_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h11));
    _zz_rob_17_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h11));
    _zz_rob_17_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h11));
    _zz_rob_17_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h11));
    _zz_rob_17_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h11));
  end

  always @(*) begin
    _zz_rob_17_isComplete_1[0] = ((head_0 == 5'h11) && retireMask[0]);
    _zz_rob_17_isComplete_1[1] = ((head_1 == 5'h11) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_18_valid[0] = ((tail_0 == 5'h12) && io_dispatch_allowMask[0]);
    _zz_rob_18_valid[1] = ((tail_1 == 5'h12) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_18_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h12));
    _zz_rob_18_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h12));
    _zz_rob_18_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h12));
    _zz_rob_18_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h12));
    _zz_rob_18_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h12));
  end

  always @(*) begin
    _zz_rob_18_isComplete_1[0] = ((head_0 == 5'h12) && retireMask[0]);
    _zz_rob_18_isComplete_1[1] = ((head_1 == 5'h12) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_19_valid[0] = ((tail_0 == 5'h13) && io_dispatch_allowMask[0]);
    _zz_rob_19_valid[1] = ((tail_1 == 5'h13) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_19_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h13));
    _zz_rob_19_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h13));
    _zz_rob_19_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h13));
    _zz_rob_19_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h13));
    _zz_rob_19_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h13));
  end

  always @(*) begin
    _zz_rob_19_isComplete_1[0] = ((head_0 == 5'h13) && retireMask[0]);
    _zz_rob_19_isComplete_1[1] = ((head_1 == 5'h13) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_20_valid[0] = ((tail_0 == 5'h14) && io_dispatch_allowMask[0]);
    _zz_rob_20_valid[1] = ((tail_1 == 5'h14) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_20_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h14));
    _zz_rob_20_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h14));
    _zz_rob_20_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h14));
    _zz_rob_20_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h14));
    _zz_rob_20_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h14));
  end

  always @(*) begin
    _zz_rob_20_isComplete_1[0] = ((head_0 == 5'h14) && retireMask[0]);
    _zz_rob_20_isComplete_1[1] = ((head_1 == 5'h14) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_21_valid[0] = ((tail_0 == 5'h15) && io_dispatch_allowMask[0]);
    _zz_rob_21_valid[1] = ((tail_1 == 5'h15) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_21_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h15));
    _zz_rob_21_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h15));
    _zz_rob_21_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h15));
    _zz_rob_21_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h15));
    _zz_rob_21_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h15));
  end

  always @(*) begin
    _zz_rob_21_isComplete_1[0] = ((head_0 == 5'h15) && retireMask[0]);
    _zz_rob_21_isComplete_1[1] = ((head_1 == 5'h15) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_22_valid[0] = ((tail_0 == 5'h16) && io_dispatch_allowMask[0]);
    _zz_rob_22_valid[1] = ((tail_1 == 5'h16) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_22_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h16));
    _zz_rob_22_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h16));
    _zz_rob_22_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h16));
    _zz_rob_22_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h16));
    _zz_rob_22_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h16));
  end

  always @(*) begin
    _zz_rob_22_isComplete_1[0] = ((head_0 == 5'h16) && retireMask[0]);
    _zz_rob_22_isComplete_1[1] = ((head_1 == 5'h16) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_23_valid[0] = ((tail_0 == 5'h17) && io_dispatch_allowMask[0]);
    _zz_rob_23_valid[1] = ((tail_1 == 5'h17) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_23_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h17));
    _zz_rob_23_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h17));
    _zz_rob_23_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h17));
    _zz_rob_23_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h17));
    _zz_rob_23_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h17));
  end

  always @(*) begin
    _zz_rob_23_isComplete_1[0] = ((head_0 == 5'h17) && retireMask[0]);
    _zz_rob_23_isComplete_1[1] = ((head_1 == 5'h17) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_24_valid[0] = ((tail_0 == 5'h18) && io_dispatch_allowMask[0]);
    _zz_rob_24_valid[1] = ((tail_1 == 5'h18) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_24_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h18));
    _zz_rob_24_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h18));
    _zz_rob_24_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h18));
    _zz_rob_24_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h18));
    _zz_rob_24_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h18));
  end

  always @(*) begin
    _zz_rob_24_isComplete_1[0] = ((head_0 == 5'h18) && retireMask[0]);
    _zz_rob_24_isComplete_1[1] = ((head_1 == 5'h18) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_25_valid[0] = ((tail_0 == 5'h19) && io_dispatch_allowMask[0]);
    _zz_rob_25_valid[1] = ((tail_1 == 5'h19) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_25_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h19));
    _zz_rob_25_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h19));
    _zz_rob_25_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h19));
    _zz_rob_25_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h19));
    _zz_rob_25_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h19));
  end

  always @(*) begin
    _zz_rob_25_isComplete_1[0] = ((head_0 == 5'h19) && retireMask[0]);
    _zz_rob_25_isComplete_1[1] = ((head_1 == 5'h19) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_26_valid[0] = ((tail_0 == 5'h1a) && io_dispatch_allowMask[0]);
    _zz_rob_26_valid[1] = ((tail_1 == 5'h1a) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_26_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h1a));
    _zz_rob_26_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h1a));
    _zz_rob_26_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h1a));
    _zz_rob_26_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h1a));
    _zz_rob_26_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h1a));
  end

  always @(*) begin
    _zz_rob_26_isComplete_1[0] = ((head_0 == 5'h1a) && retireMask[0]);
    _zz_rob_26_isComplete_1[1] = ((head_1 == 5'h1a) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_27_valid[0] = ((tail_0 == 5'h1b) && io_dispatch_allowMask[0]);
    _zz_rob_27_valid[1] = ((tail_1 == 5'h1b) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_27_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h1b));
    _zz_rob_27_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h1b));
    _zz_rob_27_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h1b));
    _zz_rob_27_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h1b));
    _zz_rob_27_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h1b));
  end

  always @(*) begin
    _zz_rob_27_isComplete_1[0] = ((head_0 == 5'h1b) && retireMask[0]);
    _zz_rob_27_isComplete_1[1] = ((head_1 == 5'h1b) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_28_valid[0] = ((tail_0 == 5'h1c) && io_dispatch_allowMask[0]);
    _zz_rob_28_valid[1] = ((tail_1 == 5'h1c) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_28_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h1c));
    _zz_rob_28_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h1c));
    _zz_rob_28_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h1c));
    _zz_rob_28_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h1c));
    _zz_rob_28_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h1c));
  end

  always @(*) begin
    _zz_rob_28_isComplete_1[0] = ((head_0 == 5'h1c) && retireMask[0]);
    _zz_rob_28_isComplete_1[1] = ((head_1 == 5'h1c) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_29_valid[0] = ((tail_0 == 5'h1d) && io_dispatch_allowMask[0]);
    _zz_rob_29_valid[1] = ((tail_1 == 5'h1d) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_29_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h1d));
    _zz_rob_29_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h1d));
    _zz_rob_29_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h1d));
    _zz_rob_29_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h1d));
    _zz_rob_29_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h1d));
  end

  always @(*) begin
    _zz_rob_29_isComplete_1[0] = ((head_0 == 5'h1d) && retireMask[0]);
    _zz_rob_29_isComplete_1[1] = ((head_1 == 5'h1d) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_30_valid[0] = ((tail_0 == 5'h1e) && io_dispatch_allowMask[0]);
    _zz_rob_30_valid[1] = ((tail_1 == 5'h1e) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_30_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h1e));
    _zz_rob_30_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h1e));
    _zz_rob_30_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h1e));
    _zz_rob_30_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h1e));
    _zz_rob_30_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h1e));
  end

  always @(*) begin
    _zz_rob_30_isComplete_1[0] = ((head_0 == 5'h1e) && retireMask[0]);
    _zz_rob_30_isComplete_1[1] = ((head_1 == 5'h1e) && retireMask[1]);
  end

  always @(*) begin
    _zz_rob_31_valid[0] = ((tail_0 == 5'h1f) && io_dispatch_allowMask[0]);
    _zz_rob_31_valid[1] = ((tail_1 == 5'h1f) && io_dispatch_allowMask[1]);
  end

  always @(*) begin
    _zz_rob_31_isComplete[0] = (io_commit_0_valid && (io_commit_0_robIdx == 5'h1f));
    _zz_rob_31_isComplete[1] = (io_commit_1_valid && (io_commit_1_robIdx == 5'h1f));
    _zz_rob_31_isComplete[2] = (io_commit_2_valid && (io_commit_2_robIdx == 5'h1f));
    _zz_rob_31_isComplete[3] = (io_commit_3_valid && (io_commit_3_robIdx == 5'h1f));
    _zz_rob_31_isComplete[4] = (io_commit_4_valid && (io_commit_4_robIdx == 5'h1f));
  end

  always @(*) begin
    _zz_rob_31_isComplete_1[0] = ((head_0 == 5'h1f) && retireMask[0]);
    _zz_rob_31_isComplete_1[1] = ((head_1 == 5'h1f) && retireMask[1]);
  end

  assign when_ROB_l76 = io_dispatch_allowMask[0];
  assign _zz_1 = ({31'd0,1'b1} <<< tail_0);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = _zz_1[4];
  assign _zz_7 = _zz_1[5];
  assign _zz_8 = _zz_1[6];
  assign _zz_9 = _zz_1[7];
  assign _zz_10 = _zz_1[8];
  assign _zz_11 = _zz_1[9];
  assign _zz_12 = _zz_1[10];
  assign _zz_13 = _zz_1[11];
  assign _zz_14 = _zz_1[12];
  assign _zz_15 = _zz_1[13];
  assign _zz_16 = _zz_1[14];
  assign _zz_17 = _zz_1[15];
  assign _zz_18 = _zz_1[16];
  assign _zz_19 = _zz_1[17];
  assign _zz_20 = _zz_1[18];
  assign _zz_21 = _zz_1[19];
  assign _zz_22 = _zz_1[20];
  assign _zz_23 = _zz_1[21];
  assign _zz_24 = _zz_1[22];
  assign _zz_25 = _zz_1[23];
  assign _zz_26 = _zz_1[24];
  assign _zz_27 = _zz_1[25];
  assign _zz_28 = _zz_1[26];
  assign _zz_29 = _zz_1[27];
  assign _zz_30 = _zz_1[28];
  assign _zz_31 = _zz_1[29];
  assign _zz_32 = _zz_1[30];
  assign _zz_33 = _zz_1[31];
  assign when_ROB_l76_1 = io_dispatch_allowMask[1];
  assign _zz_34 = ({31'd0,1'b1} <<< tail_1);
  assign _zz_35 = _zz_34[0];
  assign _zz_36 = _zz_34[1];
  assign _zz_37 = _zz_34[2];
  assign _zz_38 = _zz_34[3];
  assign _zz_39 = _zz_34[4];
  assign _zz_40 = _zz_34[5];
  assign _zz_41 = _zz_34[6];
  assign _zz_42 = _zz_34[7];
  assign _zz_43 = _zz_34[8];
  assign _zz_44 = _zz_34[9];
  assign _zz_45 = _zz_34[10];
  assign _zz_46 = _zz_34[11];
  assign _zz_47 = _zz_34[12];
  assign _zz_48 = _zz_34[13];
  assign _zz_49 = _zz_34[14];
  assign _zz_50 = _zz_34[15];
  assign _zz_51 = _zz_34[16];
  assign _zz_52 = _zz_34[17];
  assign _zz_53 = _zz_34[18];
  assign _zz_54 = _zz_34[19];
  assign _zz_55 = _zz_34[20];
  assign _zz_56 = _zz_34[21];
  assign _zz_57 = _zz_34[22];
  assign _zz_58 = _zz_34[23];
  assign _zz_59 = _zz_34[24];
  assign _zz_60 = _zz_34[25];
  assign _zz_61 = _zz_34[26];
  assign _zz_62 = _zz_34[27];
  assign _zz_63 = _zz_34[28];
  assign _zz_64 = _zz_34[29];
  assign _zz_65 = _zz_34[30];
  assign _zz_66 = _zz_34[31];
  assign _zz_67 = ({31'd0,1'b1} <<< io_commit_0_robIdx);
  assign _zz_68 = _zz_67[0];
  assign _zz_69 = _zz_67[1];
  assign _zz_70 = _zz_67[2];
  assign _zz_71 = _zz_67[3];
  assign _zz_72 = _zz_67[4];
  assign _zz_73 = _zz_67[5];
  assign _zz_74 = _zz_67[6];
  assign _zz_75 = _zz_67[7];
  assign _zz_76 = _zz_67[8];
  assign _zz_77 = _zz_67[9];
  assign _zz_78 = _zz_67[10];
  assign _zz_79 = _zz_67[11];
  assign _zz_80 = _zz_67[12];
  assign _zz_81 = _zz_67[13];
  assign _zz_82 = _zz_67[14];
  assign _zz_83 = _zz_67[15];
  assign _zz_84 = _zz_67[16];
  assign _zz_85 = _zz_67[17];
  assign _zz_86 = _zz_67[18];
  assign _zz_87 = _zz_67[19];
  assign _zz_88 = _zz_67[20];
  assign _zz_89 = _zz_67[21];
  assign _zz_90 = _zz_67[22];
  assign _zz_91 = _zz_67[23];
  assign _zz_92 = _zz_67[24];
  assign _zz_93 = _zz_67[25];
  assign _zz_94 = _zz_67[26];
  assign _zz_95 = _zz_67[27];
  assign _zz_96 = _zz_67[28];
  assign _zz_97 = _zz_67[29];
  assign _zz_98 = _zz_67[30];
  assign _zz_99 = _zz_67[31];
  assign _zz_100 = ({31'd0,1'b1} <<< io_commit_0_robIdx);
  assign _zz_101 = _zz_100[0];
  assign _zz_102 = _zz_100[1];
  assign _zz_103 = _zz_100[2];
  assign _zz_104 = _zz_100[3];
  assign _zz_105 = _zz_100[4];
  assign _zz_106 = _zz_100[5];
  assign _zz_107 = _zz_100[6];
  assign _zz_108 = _zz_100[7];
  assign _zz_109 = _zz_100[8];
  assign _zz_110 = _zz_100[9];
  assign _zz_111 = _zz_100[10];
  assign _zz_112 = _zz_100[11];
  assign _zz_113 = _zz_100[12];
  assign _zz_114 = _zz_100[13];
  assign _zz_115 = _zz_100[14];
  assign _zz_116 = _zz_100[15];
  assign _zz_117 = _zz_100[16];
  assign _zz_118 = _zz_100[17];
  assign _zz_119 = _zz_100[18];
  assign _zz_120 = _zz_100[19];
  assign _zz_121 = _zz_100[20];
  assign _zz_122 = _zz_100[21];
  assign _zz_123 = _zz_100[22];
  assign _zz_124 = _zz_100[23];
  assign _zz_125 = _zz_100[24];
  assign _zz_126 = _zz_100[25];
  assign _zz_127 = _zz_100[26];
  assign _zz_128 = _zz_100[27];
  assign _zz_129 = _zz_100[28];
  assign _zz_130 = _zz_100[29];
  assign _zz_131 = _zz_100[30];
  assign _zz_132 = _zz_100[31];
  assign _zz_io_commitROBEntries_0_pc = io_commit_0_robIdx;
  assign _zz_io_commitROBEntries_0_specialOp = _zz__zz_io_commitROBEntries_0_specialOp;
  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_pc = _zz_io_commitROBEntries_0_pc_1;
    end else begin
      io_commitROBEntries_0_pc = 32'h00000000;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_ard = _zz_io_commitROBEntries_0_ard;
    end else begin
      io_commitROBEntries_0_ard = 5'h00;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_prd = _zz_io_commitROBEntries_0_prd;
    end else begin
      io_commitROBEntries_0_prd = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_pprd = _zz_io_commitROBEntries_0_pprd;
    end else begin
      io_commitROBEntries_0_pprd = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_specialOp = _zz_io_commitROBEntries_0_specialOp;
    end else begin
      io_commitROBEntries_0_specialOp = ROBSpecialOp_nop;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_isComplete = _zz_io_commitROBEntries_0_isComplete;
    end else begin
      io_commitROBEntries_0_isComplete = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_branchResult_targetPC = _zz_io_commitROBEntries_0_branchResult_targetPC;
    end else begin
      io_commitROBEntries_0_branchResult_targetPC = 32'h00000000;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_branchResult_branchResult = _zz_io_commitROBEntries_0_branchResult_branchResult;
    end else begin
      io_commitROBEntries_0_branchResult_branchResult = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_branchResult_predictFail = _zz_io_commitROBEntries_0_branchResult_predictFail;
    end else begin
      io_commitROBEntries_0_branchResult_predictFail = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_exceptionInfo_exception = _zz_io_commitROBEntries_0_exceptionInfo_exception;
    end else begin
      io_commitROBEntries_0_exceptionInfo_exception = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_exceptionInfo_eCode = _zz_io_commitROBEntries_0_exceptionInfo_eCode;
    end else begin
      io_commitROBEntries_0_exceptionInfo_eCode = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_exceptionInfo_eSubCode = _zz_io_commitROBEntries_0_exceptionInfo_eSubCode;
    end else begin
      io_commitROBEntries_0_exceptionInfo_eSubCode = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_0_valid) begin
      io_commitROBEntries_0_valid = _zz_io_commitROBEntries_0_valid;
    end else begin
      io_commitROBEntries_0_valid = 1'b0;
    end
  end

  assign _zz_133 = ({31'd0,1'b1} <<< io_commit_1_robIdx);
  assign _zz_134 = _zz_133[0];
  assign _zz_135 = _zz_133[1];
  assign _zz_136 = _zz_133[2];
  assign _zz_137 = _zz_133[3];
  assign _zz_138 = _zz_133[4];
  assign _zz_139 = _zz_133[5];
  assign _zz_140 = _zz_133[6];
  assign _zz_141 = _zz_133[7];
  assign _zz_142 = _zz_133[8];
  assign _zz_143 = _zz_133[9];
  assign _zz_144 = _zz_133[10];
  assign _zz_145 = _zz_133[11];
  assign _zz_146 = _zz_133[12];
  assign _zz_147 = _zz_133[13];
  assign _zz_148 = _zz_133[14];
  assign _zz_149 = _zz_133[15];
  assign _zz_150 = _zz_133[16];
  assign _zz_151 = _zz_133[17];
  assign _zz_152 = _zz_133[18];
  assign _zz_153 = _zz_133[19];
  assign _zz_154 = _zz_133[20];
  assign _zz_155 = _zz_133[21];
  assign _zz_156 = _zz_133[22];
  assign _zz_157 = _zz_133[23];
  assign _zz_158 = _zz_133[24];
  assign _zz_159 = _zz_133[25];
  assign _zz_160 = _zz_133[26];
  assign _zz_161 = _zz_133[27];
  assign _zz_162 = _zz_133[28];
  assign _zz_163 = _zz_133[29];
  assign _zz_164 = _zz_133[30];
  assign _zz_165 = _zz_133[31];
  assign _zz_166 = ({31'd0,1'b1} <<< io_commit_1_robIdx);
  assign _zz_167 = _zz_166[0];
  assign _zz_168 = _zz_166[1];
  assign _zz_169 = _zz_166[2];
  assign _zz_170 = _zz_166[3];
  assign _zz_171 = _zz_166[4];
  assign _zz_172 = _zz_166[5];
  assign _zz_173 = _zz_166[6];
  assign _zz_174 = _zz_166[7];
  assign _zz_175 = _zz_166[8];
  assign _zz_176 = _zz_166[9];
  assign _zz_177 = _zz_166[10];
  assign _zz_178 = _zz_166[11];
  assign _zz_179 = _zz_166[12];
  assign _zz_180 = _zz_166[13];
  assign _zz_181 = _zz_166[14];
  assign _zz_182 = _zz_166[15];
  assign _zz_183 = _zz_166[16];
  assign _zz_184 = _zz_166[17];
  assign _zz_185 = _zz_166[18];
  assign _zz_186 = _zz_166[19];
  assign _zz_187 = _zz_166[20];
  assign _zz_188 = _zz_166[21];
  assign _zz_189 = _zz_166[22];
  assign _zz_190 = _zz_166[23];
  assign _zz_191 = _zz_166[24];
  assign _zz_192 = _zz_166[25];
  assign _zz_193 = _zz_166[26];
  assign _zz_194 = _zz_166[27];
  assign _zz_195 = _zz_166[28];
  assign _zz_196 = _zz_166[29];
  assign _zz_197 = _zz_166[30];
  assign _zz_198 = _zz_166[31];
  assign _zz_io_commitROBEntries_1_pc = io_commit_1_robIdx;
  assign _zz_io_commitROBEntries_1_specialOp = _zz__zz_io_commitROBEntries_1_specialOp;
  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_pc = _zz_io_commitROBEntries_1_pc_1;
    end else begin
      io_commitROBEntries_1_pc = 32'h00000000;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_ard = _zz_io_commitROBEntries_1_ard;
    end else begin
      io_commitROBEntries_1_ard = 5'h00;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_prd = _zz_io_commitROBEntries_1_prd;
    end else begin
      io_commitROBEntries_1_prd = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_pprd = _zz_io_commitROBEntries_1_pprd;
    end else begin
      io_commitROBEntries_1_pprd = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_specialOp = _zz_io_commitROBEntries_1_specialOp;
    end else begin
      io_commitROBEntries_1_specialOp = ROBSpecialOp_nop;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_isComplete = _zz_io_commitROBEntries_1_isComplete;
    end else begin
      io_commitROBEntries_1_isComplete = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_branchResult_targetPC = _zz_io_commitROBEntries_1_branchResult_targetPC;
    end else begin
      io_commitROBEntries_1_branchResult_targetPC = 32'h00000000;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_branchResult_branchResult = _zz_io_commitROBEntries_1_branchResult_branchResult;
    end else begin
      io_commitROBEntries_1_branchResult_branchResult = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_branchResult_predictFail = _zz_io_commitROBEntries_1_branchResult_predictFail;
    end else begin
      io_commitROBEntries_1_branchResult_predictFail = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_exceptionInfo_exception = _zz_io_commitROBEntries_1_exceptionInfo_exception;
    end else begin
      io_commitROBEntries_1_exceptionInfo_exception = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_exceptionInfo_eCode = _zz_io_commitROBEntries_1_exceptionInfo_eCode;
    end else begin
      io_commitROBEntries_1_exceptionInfo_eCode = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_exceptionInfo_eSubCode = _zz_io_commitROBEntries_1_exceptionInfo_eSubCode;
    end else begin
      io_commitROBEntries_1_exceptionInfo_eSubCode = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_1_valid) begin
      io_commitROBEntries_1_valid = _zz_io_commitROBEntries_1_valid;
    end else begin
      io_commitROBEntries_1_valid = 1'b0;
    end
  end

  assign _zz_199 = ({31'd0,1'b1} <<< io_commit_2_robIdx);
  assign _zz_200 = _zz_199[0];
  assign _zz_201 = _zz_199[1];
  assign _zz_202 = _zz_199[2];
  assign _zz_203 = _zz_199[3];
  assign _zz_204 = _zz_199[4];
  assign _zz_205 = _zz_199[5];
  assign _zz_206 = _zz_199[6];
  assign _zz_207 = _zz_199[7];
  assign _zz_208 = _zz_199[8];
  assign _zz_209 = _zz_199[9];
  assign _zz_210 = _zz_199[10];
  assign _zz_211 = _zz_199[11];
  assign _zz_212 = _zz_199[12];
  assign _zz_213 = _zz_199[13];
  assign _zz_214 = _zz_199[14];
  assign _zz_215 = _zz_199[15];
  assign _zz_216 = _zz_199[16];
  assign _zz_217 = _zz_199[17];
  assign _zz_218 = _zz_199[18];
  assign _zz_219 = _zz_199[19];
  assign _zz_220 = _zz_199[20];
  assign _zz_221 = _zz_199[21];
  assign _zz_222 = _zz_199[22];
  assign _zz_223 = _zz_199[23];
  assign _zz_224 = _zz_199[24];
  assign _zz_225 = _zz_199[25];
  assign _zz_226 = _zz_199[26];
  assign _zz_227 = _zz_199[27];
  assign _zz_228 = _zz_199[28];
  assign _zz_229 = _zz_199[29];
  assign _zz_230 = _zz_199[30];
  assign _zz_231 = _zz_199[31];
  assign _zz_232 = ({31'd0,1'b1} <<< io_commit_2_robIdx);
  assign _zz_233 = _zz_232[0];
  assign _zz_234 = _zz_232[1];
  assign _zz_235 = _zz_232[2];
  assign _zz_236 = _zz_232[3];
  assign _zz_237 = _zz_232[4];
  assign _zz_238 = _zz_232[5];
  assign _zz_239 = _zz_232[6];
  assign _zz_240 = _zz_232[7];
  assign _zz_241 = _zz_232[8];
  assign _zz_242 = _zz_232[9];
  assign _zz_243 = _zz_232[10];
  assign _zz_244 = _zz_232[11];
  assign _zz_245 = _zz_232[12];
  assign _zz_246 = _zz_232[13];
  assign _zz_247 = _zz_232[14];
  assign _zz_248 = _zz_232[15];
  assign _zz_249 = _zz_232[16];
  assign _zz_250 = _zz_232[17];
  assign _zz_251 = _zz_232[18];
  assign _zz_252 = _zz_232[19];
  assign _zz_253 = _zz_232[20];
  assign _zz_254 = _zz_232[21];
  assign _zz_255 = _zz_232[22];
  assign _zz_256 = _zz_232[23];
  assign _zz_257 = _zz_232[24];
  assign _zz_258 = _zz_232[25];
  assign _zz_259 = _zz_232[26];
  assign _zz_260 = _zz_232[27];
  assign _zz_261 = _zz_232[28];
  assign _zz_262 = _zz_232[29];
  assign _zz_263 = _zz_232[30];
  assign _zz_264 = _zz_232[31];
  assign _zz_io_commitROBEntries_2_pc = io_commit_2_robIdx;
  assign _zz_io_commitROBEntries_2_specialOp = _zz__zz_io_commitROBEntries_2_specialOp;
  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_pc = _zz_io_commitROBEntries_2_pc_1;
    end else begin
      io_commitROBEntries_2_pc = 32'h00000000;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_ard = _zz_io_commitROBEntries_2_ard;
    end else begin
      io_commitROBEntries_2_ard = 5'h00;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_prd = _zz_io_commitROBEntries_2_prd;
    end else begin
      io_commitROBEntries_2_prd = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_pprd = _zz_io_commitROBEntries_2_pprd;
    end else begin
      io_commitROBEntries_2_pprd = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_specialOp = _zz_io_commitROBEntries_2_specialOp;
    end else begin
      io_commitROBEntries_2_specialOp = ROBSpecialOp_nop;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_isComplete = _zz_io_commitROBEntries_2_isComplete;
    end else begin
      io_commitROBEntries_2_isComplete = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_branchResult_targetPC = _zz_io_commitROBEntries_2_branchResult_targetPC;
    end else begin
      io_commitROBEntries_2_branchResult_targetPC = 32'h00000000;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_branchResult_branchResult = _zz_io_commitROBEntries_2_branchResult_branchResult;
    end else begin
      io_commitROBEntries_2_branchResult_branchResult = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_branchResult_predictFail = _zz_io_commitROBEntries_2_branchResult_predictFail;
    end else begin
      io_commitROBEntries_2_branchResult_predictFail = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_exceptionInfo_exception = _zz_io_commitROBEntries_2_exceptionInfo_exception;
    end else begin
      io_commitROBEntries_2_exceptionInfo_exception = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_exceptionInfo_eCode = _zz_io_commitROBEntries_2_exceptionInfo_eCode;
    end else begin
      io_commitROBEntries_2_exceptionInfo_eCode = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_exceptionInfo_eSubCode = _zz_io_commitROBEntries_2_exceptionInfo_eSubCode;
    end else begin
      io_commitROBEntries_2_exceptionInfo_eSubCode = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_2_valid) begin
      io_commitROBEntries_2_valid = _zz_io_commitROBEntries_2_valid;
    end else begin
      io_commitROBEntries_2_valid = 1'b0;
    end
  end

  assign _zz_265 = ({31'd0,1'b1} <<< io_commit_3_robIdx);
  assign _zz_266 = _zz_265[0];
  assign _zz_267 = _zz_265[1];
  assign _zz_268 = _zz_265[2];
  assign _zz_269 = _zz_265[3];
  assign _zz_270 = _zz_265[4];
  assign _zz_271 = _zz_265[5];
  assign _zz_272 = _zz_265[6];
  assign _zz_273 = _zz_265[7];
  assign _zz_274 = _zz_265[8];
  assign _zz_275 = _zz_265[9];
  assign _zz_276 = _zz_265[10];
  assign _zz_277 = _zz_265[11];
  assign _zz_278 = _zz_265[12];
  assign _zz_279 = _zz_265[13];
  assign _zz_280 = _zz_265[14];
  assign _zz_281 = _zz_265[15];
  assign _zz_282 = _zz_265[16];
  assign _zz_283 = _zz_265[17];
  assign _zz_284 = _zz_265[18];
  assign _zz_285 = _zz_265[19];
  assign _zz_286 = _zz_265[20];
  assign _zz_287 = _zz_265[21];
  assign _zz_288 = _zz_265[22];
  assign _zz_289 = _zz_265[23];
  assign _zz_290 = _zz_265[24];
  assign _zz_291 = _zz_265[25];
  assign _zz_292 = _zz_265[26];
  assign _zz_293 = _zz_265[27];
  assign _zz_294 = _zz_265[28];
  assign _zz_295 = _zz_265[29];
  assign _zz_296 = _zz_265[30];
  assign _zz_297 = _zz_265[31];
  assign _zz_298 = ({31'd0,1'b1} <<< io_commit_3_robIdx);
  assign _zz_299 = _zz_298[0];
  assign _zz_300 = _zz_298[1];
  assign _zz_301 = _zz_298[2];
  assign _zz_302 = _zz_298[3];
  assign _zz_303 = _zz_298[4];
  assign _zz_304 = _zz_298[5];
  assign _zz_305 = _zz_298[6];
  assign _zz_306 = _zz_298[7];
  assign _zz_307 = _zz_298[8];
  assign _zz_308 = _zz_298[9];
  assign _zz_309 = _zz_298[10];
  assign _zz_310 = _zz_298[11];
  assign _zz_311 = _zz_298[12];
  assign _zz_312 = _zz_298[13];
  assign _zz_313 = _zz_298[14];
  assign _zz_314 = _zz_298[15];
  assign _zz_315 = _zz_298[16];
  assign _zz_316 = _zz_298[17];
  assign _zz_317 = _zz_298[18];
  assign _zz_318 = _zz_298[19];
  assign _zz_319 = _zz_298[20];
  assign _zz_320 = _zz_298[21];
  assign _zz_321 = _zz_298[22];
  assign _zz_322 = _zz_298[23];
  assign _zz_323 = _zz_298[24];
  assign _zz_324 = _zz_298[25];
  assign _zz_325 = _zz_298[26];
  assign _zz_326 = _zz_298[27];
  assign _zz_327 = _zz_298[28];
  assign _zz_328 = _zz_298[29];
  assign _zz_329 = _zz_298[30];
  assign _zz_330 = _zz_298[31];
  assign _zz_io_commitROBEntries_3_pc = io_commit_3_robIdx;
  assign _zz_io_commitROBEntries_3_specialOp = _zz__zz_io_commitROBEntries_3_specialOp;
  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_pc = _zz_io_commitROBEntries_3_pc_1;
    end else begin
      io_commitROBEntries_3_pc = 32'h00000000;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_ard = _zz_io_commitROBEntries_3_ard;
    end else begin
      io_commitROBEntries_3_ard = 5'h00;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_prd = _zz_io_commitROBEntries_3_prd;
    end else begin
      io_commitROBEntries_3_prd = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_pprd = _zz_io_commitROBEntries_3_pprd;
    end else begin
      io_commitROBEntries_3_pprd = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_specialOp = _zz_io_commitROBEntries_3_specialOp;
    end else begin
      io_commitROBEntries_3_specialOp = ROBSpecialOp_nop;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_isComplete = _zz_io_commitROBEntries_3_isComplete;
    end else begin
      io_commitROBEntries_3_isComplete = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_branchResult_targetPC = _zz_io_commitROBEntries_3_branchResult_targetPC;
    end else begin
      io_commitROBEntries_3_branchResult_targetPC = 32'h00000000;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_branchResult_branchResult = _zz_io_commitROBEntries_3_branchResult_branchResult;
    end else begin
      io_commitROBEntries_3_branchResult_branchResult = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_branchResult_predictFail = _zz_io_commitROBEntries_3_branchResult_predictFail;
    end else begin
      io_commitROBEntries_3_branchResult_predictFail = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_exceptionInfo_exception = _zz_io_commitROBEntries_3_exceptionInfo_exception;
    end else begin
      io_commitROBEntries_3_exceptionInfo_exception = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_exceptionInfo_eCode = _zz_io_commitROBEntries_3_exceptionInfo_eCode;
    end else begin
      io_commitROBEntries_3_exceptionInfo_eCode = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_exceptionInfo_eSubCode = _zz_io_commitROBEntries_3_exceptionInfo_eSubCode;
    end else begin
      io_commitROBEntries_3_exceptionInfo_eSubCode = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_3_valid) begin
      io_commitROBEntries_3_valid = _zz_io_commitROBEntries_3_valid;
    end else begin
      io_commitROBEntries_3_valid = 1'b0;
    end
  end

  assign _zz_331 = ({31'd0,1'b1} <<< io_commit_4_robIdx);
  assign _zz_332 = _zz_331[0];
  assign _zz_333 = _zz_331[1];
  assign _zz_334 = _zz_331[2];
  assign _zz_335 = _zz_331[3];
  assign _zz_336 = _zz_331[4];
  assign _zz_337 = _zz_331[5];
  assign _zz_338 = _zz_331[6];
  assign _zz_339 = _zz_331[7];
  assign _zz_340 = _zz_331[8];
  assign _zz_341 = _zz_331[9];
  assign _zz_342 = _zz_331[10];
  assign _zz_343 = _zz_331[11];
  assign _zz_344 = _zz_331[12];
  assign _zz_345 = _zz_331[13];
  assign _zz_346 = _zz_331[14];
  assign _zz_347 = _zz_331[15];
  assign _zz_348 = _zz_331[16];
  assign _zz_349 = _zz_331[17];
  assign _zz_350 = _zz_331[18];
  assign _zz_351 = _zz_331[19];
  assign _zz_352 = _zz_331[20];
  assign _zz_353 = _zz_331[21];
  assign _zz_354 = _zz_331[22];
  assign _zz_355 = _zz_331[23];
  assign _zz_356 = _zz_331[24];
  assign _zz_357 = _zz_331[25];
  assign _zz_358 = _zz_331[26];
  assign _zz_359 = _zz_331[27];
  assign _zz_360 = _zz_331[28];
  assign _zz_361 = _zz_331[29];
  assign _zz_362 = _zz_331[30];
  assign _zz_363 = _zz_331[31];
  assign _zz_364 = ({31'd0,1'b1} <<< io_commit_4_robIdx);
  assign _zz_365 = _zz_364[0];
  assign _zz_366 = _zz_364[1];
  assign _zz_367 = _zz_364[2];
  assign _zz_368 = _zz_364[3];
  assign _zz_369 = _zz_364[4];
  assign _zz_370 = _zz_364[5];
  assign _zz_371 = _zz_364[6];
  assign _zz_372 = _zz_364[7];
  assign _zz_373 = _zz_364[8];
  assign _zz_374 = _zz_364[9];
  assign _zz_375 = _zz_364[10];
  assign _zz_376 = _zz_364[11];
  assign _zz_377 = _zz_364[12];
  assign _zz_378 = _zz_364[13];
  assign _zz_379 = _zz_364[14];
  assign _zz_380 = _zz_364[15];
  assign _zz_381 = _zz_364[16];
  assign _zz_382 = _zz_364[17];
  assign _zz_383 = _zz_364[18];
  assign _zz_384 = _zz_364[19];
  assign _zz_385 = _zz_364[20];
  assign _zz_386 = _zz_364[21];
  assign _zz_387 = _zz_364[22];
  assign _zz_388 = _zz_364[23];
  assign _zz_389 = _zz_364[24];
  assign _zz_390 = _zz_364[25];
  assign _zz_391 = _zz_364[26];
  assign _zz_392 = _zz_364[27];
  assign _zz_393 = _zz_364[28];
  assign _zz_394 = _zz_364[29];
  assign _zz_395 = _zz_364[30];
  assign _zz_396 = _zz_364[31];
  assign _zz_io_commitROBEntries_4_pc = io_commit_4_robIdx;
  assign _zz_io_commitROBEntries_4_specialOp = _zz__zz_io_commitROBEntries_4_specialOp;
  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_pc = _zz_io_commitROBEntries_4_pc_1;
    end else begin
      io_commitROBEntries_4_pc = 32'h00000000;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_ard = _zz_io_commitROBEntries_4_ard;
    end else begin
      io_commitROBEntries_4_ard = 5'h00;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_prd = _zz_io_commitROBEntries_4_prd;
    end else begin
      io_commitROBEntries_4_prd = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_pprd = _zz_io_commitROBEntries_4_pprd;
    end else begin
      io_commitROBEntries_4_pprd = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_specialOp = _zz_io_commitROBEntries_4_specialOp;
    end else begin
      io_commitROBEntries_4_specialOp = ROBSpecialOp_nop;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_isComplete = _zz_io_commitROBEntries_4_isComplete;
    end else begin
      io_commitROBEntries_4_isComplete = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_branchResult_targetPC = _zz_io_commitROBEntries_4_branchResult_targetPC;
    end else begin
      io_commitROBEntries_4_branchResult_targetPC = 32'h00000000;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_branchResult_branchResult = _zz_io_commitROBEntries_4_branchResult_branchResult;
    end else begin
      io_commitROBEntries_4_branchResult_branchResult = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_branchResult_predictFail = _zz_io_commitROBEntries_4_branchResult_predictFail;
    end else begin
      io_commitROBEntries_4_branchResult_predictFail = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_exceptionInfo_exception = _zz_io_commitROBEntries_4_exceptionInfo_exception;
    end else begin
      io_commitROBEntries_4_exceptionInfo_exception = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_exceptionInfo_eCode = _zz_io_commitROBEntries_4_exceptionInfo_eCode;
    end else begin
      io_commitROBEntries_4_exceptionInfo_eCode = 6'h00;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_exceptionInfo_eSubCode = _zz_io_commitROBEntries_4_exceptionInfo_eSubCode;
    end else begin
      io_commitROBEntries_4_exceptionInfo_eSubCode = 1'b0;
    end
  end

  always @(*) begin
    if(io_commit_4_valid) begin
      io_commitROBEntries_4_valid = _zz_io_commitROBEntries_4_valid;
    end else begin
      io_commitROBEntries_4_valid = 1'b0;
    end
  end

  always @(*) begin
    inhibitNextRetireMask[0] = (((((_zz_stage_updateBPU_0_isJumpInst == ROBSpecialOp_lsuAction) || (_zz_stage_updateBPU_0_isJumpInst == ROBSpecialOp_ll)) || (_zz_stage_updateBPU_0_isJumpInst == ROBSpecialOp_writeCSR)) || (_zz_stage_updateBPU_0_isJumpInst == ROBSpecialOp_ertn)) || _zz_stage_updateBPU_0_predictFail);
    inhibitNextRetireMask[1] = (((((_zz_stage_updateBPU_1_isJumpInst == ROBSpecialOp_lsuAction) || (_zz_stage_updateBPU_1_isJumpInst == ROBSpecialOp_ll)) || (_zz_stage_updateBPU_1_isJumpInst == ROBSpecialOp_writeCSR)) || (_zz_stage_updateBPU_1_isJumpInst == ROBSpecialOp_ertn)) || _zz_stage_updateBPU_1_predictFail);
  end

  assign _zz_retireEPC = flushMask[0];
  assign retireEPC = (idleEn ? retireSNPC_0 : (_zz_retireEPC ? retirePC_0 : retirePC_1));
  assign retireRealEROBIdx = (_zz_retireEPC ? retireEROBIdx_0 : retireEROBIdx_1);
  assign retireRealECode = (idleEn ? 6'h00 : (_zz_retireEPC ? retireECode_0 : retireECode_1));
  assign retireRealESubCode = (idleEn ? 1'b0 : (_zz_retireEPC ? retireESubCode_0 : retireESubCode_1));
  assign ertn = (|(ertnMask & retireMask));
  assign normalException = ((_zz_retireEPC ? normalExceptionMask[0] : normalExceptionMask[1]) || idleEn);
  assign tlbrException = (_zz_retireEPC ? tlbrExceptionMask[0] : tlbrExceptionMask[1]);
  assign falseTaken = (_zz_retireEPC ? falseTakenMask[0] : falseTakenMask[1]);
  assign snpc = (_zz_retireEPC ? retireSNPC_0 : retireSNPC_1);
  assign targetPC = (_zz_retireEPC ? retireTargetPC_0 : retireTargetPC_1);
  assign noPPRDMaskMid_0_0 = noPPRDMask[0];
  assign freePRFIdxMid_0_0 = _zz_noPPRDMask;
  assign noPPRDMaskMid_0_1 = noPPRDMask[1];
  assign freePRFIdxMid_0_1 = _zz_noPPRDMask;
  assign noPPRDMaskMid_1_0 = ((&_zz_noPPRDMaskMid_1_0[0 : 0]) ? noPPRDMaskMid_0_0 : noPPRDMaskMid_0_1);
  assign freePRFIdxMid_1_0 = ((&_zz_freePRFIdxMid_1_0[0 : 0]) ? freePRFIdxMid_0_0 : freePRFIdxMid_0_1);
  assign noPPRDMaskMid_1_1 = ((&_zz_noPPRDMaskMid_1_1[1 : 0]) ? noPPRDMaskMid_0_1 : 1'b0);
  assign freePRFIdxMid_1_1 = ((&_zz_freePRFIdxMid_1_1[1 : 0]) ? freePRFIdxMid_0_1 : 6'h00);
  assign stage_retireARAT_0_ard = _zz_stage_retireARAT_0_ard;
  assign stage_retireARAT_0_prd = _zz_stage_retireARAT_0_prd;
  assign stage_retireARAT_0_wen = retireMask[0];
  always @(*) begin
    noPPRDMask[0] = (_zz_noPPRDMask == 6'h00);
    noPPRDMask[1] = (_zz_noPPRDMask_1 == 6'h00);
  end

  always @(*) begin
    lsuActionMask[0] = (_zz_stage_updateBPU_0_isJumpInst == ROBSpecialOp_lsuAction);
    lsuActionMask[1] = (_zz_stage_updateBPU_1_isJumpInst == ROBSpecialOp_lsuAction);
  end

  always @(*) begin
    llMask[0] = (_zz_stage_updateBPU_0_isJumpInst == ROBSpecialOp_ll);
    llMask[1] = (_zz_stage_updateBPU_1_isJumpInst == ROBSpecialOp_ll);
  end

  always @(*) begin
    writeCSRMask[0] = (_zz_stage_updateBPU_0_isJumpInst == ROBSpecialOp_writeCSR);
    writeCSRMask[1] = (_zz_stage_updateBPU_1_isJumpInst == ROBSpecialOp_writeCSR);
  end

  always @(*) begin
    ertnMask[0] = (_zz_stage_updateBPU_0_isJumpInst == ROBSpecialOp_ertn);
    ertnMask[1] = (_zz_stage_updateBPU_1_isJumpInst == ROBSpecialOp_ertn);
  end

  always @(*) begin
    normalExceptionMask[0] = ((_zz_retireMask && _zz_retireMask_1) && ((_zz_normalExceptionMask != 6'h3f) || (_zz_normalExceptionMask_1 != 1'b0)));
    normalExceptionMask[1] = ((_zz_retireMask_3 && _zz_retireMask_4) && ((_zz_normalExceptionMask_2 != 6'h3f) || (_zz_normalExceptionMask_3 != 1'b0)));
  end

  always @(*) begin
    tlbrExceptionMask[0] = ((_zz_retireMask && _zz_retireMask_1) && ((_zz_normalExceptionMask == 6'h3f) && (_zz_normalExceptionMask_1 == 1'b0)));
    tlbrExceptionMask[1] = ((_zz_retireMask_3 && _zz_retireMask_4) && ((_zz_normalExceptionMask_2 == 6'h3f) && (_zz_normalExceptionMask_3 == 1'b0)));
  end

  always @(*) begin
    falseTakenMask[0] = ((_zz_retireMask && (! _zz_stage_updateBPU_0_taken)) && _zz_stage_updateBPU_0_predictFail);
    falseTakenMask[1] = ((_zz_retireMask_3 && (! _zz_stage_updateBPU_1_taken)) && _zz_stage_updateBPU_1_predictFail);
  end

  assign retirePC_0 = _zz_retirePC_0;
  assign retireEROBIdx_0 = head_0;
  assign retireECode_0 = _zz_normalExceptionMask;
  assign retireESubCode_0 = _zz_normalExceptionMask_1;
  assign retireSNPC_0 = (_zz_retirePC_0 + 32'h00000004);
  assign retireTargetPC_0 = _zz_retireTargetPC_0;
  assign stage_freePRFIdx_0 = freePRFIdxMid_1_0;
  assign stage_retireROBIdx_0 = head_0;
  assign stage_retireEn_0 = retireMask[0];
  assign stage_updateBPU_0_pc = retirePC_0;
  assign stage_updateBPU_0_isJumpInst = (_zz_stage_updateBPU_0_isJumpInst == ROBSpecialOp_bpuUpdate);
  assign stage_updateBPU_0_taken = _zz_stage_updateBPU_0_taken;
  assign stage_updateBPU_0_predictFail = _zz_stage_updateBPU_0_predictFail;
  assign stage_updateBPU_0_target = retireTargetPC_0;
  assign stage_retireARAT_1_ard = _zz_stage_retireARAT_1_ard;
  assign stage_retireARAT_1_prd = _zz_stage_retireARAT_1_prd;
  assign stage_retireARAT_1_wen = retireMask[1];
  assign retirePC_1 = _zz_retirePC_1;
  assign retireEROBIdx_1 = head_1;
  assign retireECode_1 = _zz_normalExceptionMask_2;
  assign retireESubCode_1 = _zz_normalExceptionMask_3;
  assign retireSNPC_1 = (_zz_retirePC_1 + 32'h00000004);
  assign retireTargetPC_1 = _zz_retireTargetPC_1;
  assign stage_freePRFIdx_1 = freePRFIdxMid_1_1;
  assign stage_retireROBIdx_1 = head_1;
  assign stage_retireEn_1 = retireMask[1];
  assign stage_updateBPU_1_pc = retirePC_1;
  assign stage_updateBPU_1_isJumpInst = (_zz_stage_updateBPU_1_isJumpInst == ROBSpecialOp_bpuUpdate);
  assign stage_updateBPU_1_taken = _zz_stage_updateBPU_1_taken;
  assign stage_updateBPU_1_predictFail = _zz_stage_updateBPU_1_predictFail;
  assign stage_updateBPU_1_target = retireTargetPC_1;
  assign _zz_stage_freePRFNum = ((~ noPPRDMask) & retireMask);
  assign stage_freePRFNum = _zz_stage_freePRFNum_1;
  assign stage_wakeupMem = (|(lsuActionMask & retireMask));
  assign stage_retireLLBitUpdate = (|(llMask & retireMask));
  assign stage_retireWriteCSR = (|(writeCSRMask & retireMask));
  assign stage_retireERTN = ertn;
  assign stage_retireNormalException = normalException;
  assign stage_retireTLBRException = tlbrException;
  assign stage_retireEPC = retireEPC;
  assign stage_retireEROBIdx = retireRealEROBIdx;
  assign stage_retireECode = retireRealECode;
  assign stage_retireESubCode = retireRealESubCode;
  assign stage_flush = flush;
  assign stage_redirectPC = (normalException ? io_csrCtrl_eentry : (tlbrException ? io_csrCtrl_tlbrentry : (ertn ? io_csrCtrl_era : (falseTaken ? snpc : targetPC))));
  assign io_dispatch_availMask = stageReg_availROBMask;
  assign io_retireARAT_0_ard = stageReg_retireARAT_0_ard;
  assign io_retireARAT_0_prd = stageReg_retireARAT_0_prd;
  assign io_retireARAT_0_wen = stageReg_retireARAT_0_wen;
  assign io_retireARAT_1_ard = stageReg_retireARAT_1_ard;
  assign io_retireARAT_1_prd = stageReg_retireARAT_1_prd;
  assign io_retireARAT_1_wen = stageReg_retireARAT_1_wen;
  assign io_retireFreeList_prfIdx_0 = stageReg_freePRFIdx_0;
  assign io_retireFreeList_prfIdx_1 = stageReg_freePRFIdx_1;
  assign io_retireFreeList_writeNum = stageReg_freePRFNum;
  assign io_retireFreeList_delayedFlush = delayedFlush;
  assign io_retireLSU_robIdx_0 = stageReg_retireROBIdx_0;
  assign io_retireLSU_robIdx_1 = stageReg_retireROBIdx_1;
  assign io_retireLSU_allowRetire_0 = stageReg_retireEn_0;
  assign io_retireLSU_allowRetire_1 = stageReg_retireEn_1;
  assign io_wakeupMem = stageReg_wakeupMem;
  assign io_csrCtrl_llBitUpdate = stageReg_retireLLBitUpdate;
  assign io_csrCtrl_writeCSR = stageReg_retireWriteCSR;
  assign io_csrCtrl_ertn = stageReg_retireERTN;
  assign io_csrCtrl_normalException = stageReg_retireNormalException;
  assign io_csrCtrl_tlbrException = stageReg_retireTLBRException;
  assign io_csrCtrl_epc = stageReg_retireEPC;
  assign io_csrCtrl_eROBIdx = stageReg_retireEROBIdx;
  assign io_csrCtrl_eCode = stageReg_retireECode;
  assign io_csrCtrl_eSubCode = stageReg_retireESubCode;
  assign io_flush = stageReg_flush;
  assign io_redirectPC = stageReg_redirectPC;
  assign io_updateBPU_0_valid = stageReg_retireEn_0;
  assign io_updateBPU_0_payload_pc = stageReg_updateBPU_0_pc;
  assign io_updateBPU_0_payload_isJumpInst = stageReg_updateBPU_0_isJumpInst;
  assign io_updateBPU_0_payload_taken = stageReg_updateBPU_0_taken;
  assign io_updateBPU_0_payload_predictFail = stageReg_updateBPU_0_predictFail;
  assign io_updateBPU_0_payload_target = stageReg_updateBPU_0_target;
  assign io_updateBPU_1_valid = stageReg_retireEn_1;
  assign io_updateBPU_1_payload_pc = stageReg_updateBPU_1_pc;
  assign io_updateBPU_1_payload_isJumpInst = stageReg_updateBPU_1_isJumpInst;
  assign io_updateBPU_1_payload_taken = stageReg_updateBPU_1_taken;
  assign io_updateBPU_1_payload_predictFail = stageReg_updateBPU_1_predictFail;
  assign io_updateBPU_1_payload_target = stageReg_updateBPU_1_target;
  always @(posedge aclk) begin
    if(!aresetn) begin
      rob_0_pc <= 32'h00000000;
      rob_0_ard <= 5'h00;
      rob_0_prd <= 6'h00;
      rob_0_pprd <= 6'h00;
      rob_0_specialOp <= ROBSpecialOp_nop;
      rob_0_isComplete <= 1'b0;
      rob_0_branchResult_targetPC <= 32'h00000000;
      rob_0_branchResult_branchResult <= 1'b0;
      rob_0_branchResult_predictFail <= 1'b0;
      rob_0_exceptionInfo_exception <= 1'b0;
      rob_0_exceptionInfo_eCode <= 6'h00;
      rob_0_exceptionInfo_eSubCode <= 1'b0;
      rob_0_valid <= 1'b0;
      rob_1_pc <= 32'h00000000;
      rob_1_ard <= 5'h00;
      rob_1_prd <= 6'h00;
      rob_1_pprd <= 6'h00;
      rob_1_specialOp <= ROBSpecialOp_nop;
      rob_1_isComplete <= 1'b0;
      rob_1_branchResult_targetPC <= 32'h00000000;
      rob_1_branchResult_branchResult <= 1'b0;
      rob_1_branchResult_predictFail <= 1'b0;
      rob_1_exceptionInfo_exception <= 1'b0;
      rob_1_exceptionInfo_eCode <= 6'h00;
      rob_1_exceptionInfo_eSubCode <= 1'b0;
      rob_1_valid <= 1'b0;
      rob_2_pc <= 32'h00000000;
      rob_2_ard <= 5'h00;
      rob_2_prd <= 6'h00;
      rob_2_pprd <= 6'h00;
      rob_2_specialOp <= ROBSpecialOp_nop;
      rob_2_isComplete <= 1'b0;
      rob_2_branchResult_targetPC <= 32'h00000000;
      rob_2_branchResult_branchResult <= 1'b0;
      rob_2_branchResult_predictFail <= 1'b0;
      rob_2_exceptionInfo_exception <= 1'b0;
      rob_2_exceptionInfo_eCode <= 6'h00;
      rob_2_exceptionInfo_eSubCode <= 1'b0;
      rob_2_valid <= 1'b0;
      rob_3_pc <= 32'h00000000;
      rob_3_ard <= 5'h00;
      rob_3_prd <= 6'h00;
      rob_3_pprd <= 6'h00;
      rob_3_specialOp <= ROBSpecialOp_nop;
      rob_3_isComplete <= 1'b0;
      rob_3_branchResult_targetPC <= 32'h00000000;
      rob_3_branchResult_branchResult <= 1'b0;
      rob_3_branchResult_predictFail <= 1'b0;
      rob_3_exceptionInfo_exception <= 1'b0;
      rob_3_exceptionInfo_eCode <= 6'h00;
      rob_3_exceptionInfo_eSubCode <= 1'b0;
      rob_3_valid <= 1'b0;
      rob_4_pc <= 32'h00000000;
      rob_4_ard <= 5'h00;
      rob_4_prd <= 6'h00;
      rob_4_pprd <= 6'h00;
      rob_4_specialOp <= ROBSpecialOp_nop;
      rob_4_isComplete <= 1'b0;
      rob_4_branchResult_targetPC <= 32'h00000000;
      rob_4_branchResult_branchResult <= 1'b0;
      rob_4_branchResult_predictFail <= 1'b0;
      rob_4_exceptionInfo_exception <= 1'b0;
      rob_4_exceptionInfo_eCode <= 6'h00;
      rob_4_exceptionInfo_eSubCode <= 1'b0;
      rob_4_valid <= 1'b0;
      rob_5_pc <= 32'h00000000;
      rob_5_ard <= 5'h00;
      rob_5_prd <= 6'h00;
      rob_5_pprd <= 6'h00;
      rob_5_specialOp <= ROBSpecialOp_nop;
      rob_5_isComplete <= 1'b0;
      rob_5_branchResult_targetPC <= 32'h00000000;
      rob_5_branchResult_branchResult <= 1'b0;
      rob_5_branchResult_predictFail <= 1'b0;
      rob_5_exceptionInfo_exception <= 1'b0;
      rob_5_exceptionInfo_eCode <= 6'h00;
      rob_5_exceptionInfo_eSubCode <= 1'b0;
      rob_5_valid <= 1'b0;
      rob_6_pc <= 32'h00000000;
      rob_6_ard <= 5'h00;
      rob_6_prd <= 6'h00;
      rob_6_pprd <= 6'h00;
      rob_6_specialOp <= ROBSpecialOp_nop;
      rob_6_isComplete <= 1'b0;
      rob_6_branchResult_targetPC <= 32'h00000000;
      rob_6_branchResult_branchResult <= 1'b0;
      rob_6_branchResult_predictFail <= 1'b0;
      rob_6_exceptionInfo_exception <= 1'b0;
      rob_6_exceptionInfo_eCode <= 6'h00;
      rob_6_exceptionInfo_eSubCode <= 1'b0;
      rob_6_valid <= 1'b0;
      rob_7_pc <= 32'h00000000;
      rob_7_ard <= 5'h00;
      rob_7_prd <= 6'h00;
      rob_7_pprd <= 6'h00;
      rob_7_specialOp <= ROBSpecialOp_nop;
      rob_7_isComplete <= 1'b0;
      rob_7_branchResult_targetPC <= 32'h00000000;
      rob_7_branchResult_branchResult <= 1'b0;
      rob_7_branchResult_predictFail <= 1'b0;
      rob_7_exceptionInfo_exception <= 1'b0;
      rob_7_exceptionInfo_eCode <= 6'h00;
      rob_7_exceptionInfo_eSubCode <= 1'b0;
      rob_7_valid <= 1'b0;
      rob_8_pc <= 32'h00000000;
      rob_8_ard <= 5'h00;
      rob_8_prd <= 6'h00;
      rob_8_pprd <= 6'h00;
      rob_8_specialOp <= ROBSpecialOp_nop;
      rob_8_isComplete <= 1'b0;
      rob_8_branchResult_targetPC <= 32'h00000000;
      rob_8_branchResult_branchResult <= 1'b0;
      rob_8_branchResult_predictFail <= 1'b0;
      rob_8_exceptionInfo_exception <= 1'b0;
      rob_8_exceptionInfo_eCode <= 6'h00;
      rob_8_exceptionInfo_eSubCode <= 1'b0;
      rob_8_valid <= 1'b0;
      rob_9_pc <= 32'h00000000;
      rob_9_ard <= 5'h00;
      rob_9_prd <= 6'h00;
      rob_9_pprd <= 6'h00;
      rob_9_specialOp <= ROBSpecialOp_nop;
      rob_9_isComplete <= 1'b0;
      rob_9_branchResult_targetPC <= 32'h00000000;
      rob_9_branchResult_branchResult <= 1'b0;
      rob_9_branchResult_predictFail <= 1'b0;
      rob_9_exceptionInfo_exception <= 1'b0;
      rob_9_exceptionInfo_eCode <= 6'h00;
      rob_9_exceptionInfo_eSubCode <= 1'b0;
      rob_9_valid <= 1'b0;
      rob_10_pc <= 32'h00000000;
      rob_10_ard <= 5'h00;
      rob_10_prd <= 6'h00;
      rob_10_pprd <= 6'h00;
      rob_10_specialOp <= ROBSpecialOp_nop;
      rob_10_isComplete <= 1'b0;
      rob_10_branchResult_targetPC <= 32'h00000000;
      rob_10_branchResult_branchResult <= 1'b0;
      rob_10_branchResult_predictFail <= 1'b0;
      rob_10_exceptionInfo_exception <= 1'b0;
      rob_10_exceptionInfo_eCode <= 6'h00;
      rob_10_exceptionInfo_eSubCode <= 1'b0;
      rob_10_valid <= 1'b0;
      rob_11_pc <= 32'h00000000;
      rob_11_ard <= 5'h00;
      rob_11_prd <= 6'h00;
      rob_11_pprd <= 6'h00;
      rob_11_specialOp <= ROBSpecialOp_nop;
      rob_11_isComplete <= 1'b0;
      rob_11_branchResult_targetPC <= 32'h00000000;
      rob_11_branchResult_branchResult <= 1'b0;
      rob_11_branchResult_predictFail <= 1'b0;
      rob_11_exceptionInfo_exception <= 1'b0;
      rob_11_exceptionInfo_eCode <= 6'h00;
      rob_11_exceptionInfo_eSubCode <= 1'b0;
      rob_11_valid <= 1'b0;
      rob_12_pc <= 32'h00000000;
      rob_12_ard <= 5'h00;
      rob_12_prd <= 6'h00;
      rob_12_pprd <= 6'h00;
      rob_12_specialOp <= ROBSpecialOp_nop;
      rob_12_isComplete <= 1'b0;
      rob_12_branchResult_targetPC <= 32'h00000000;
      rob_12_branchResult_branchResult <= 1'b0;
      rob_12_branchResult_predictFail <= 1'b0;
      rob_12_exceptionInfo_exception <= 1'b0;
      rob_12_exceptionInfo_eCode <= 6'h00;
      rob_12_exceptionInfo_eSubCode <= 1'b0;
      rob_12_valid <= 1'b0;
      rob_13_pc <= 32'h00000000;
      rob_13_ard <= 5'h00;
      rob_13_prd <= 6'h00;
      rob_13_pprd <= 6'h00;
      rob_13_specialOp <= ROBSpecialOp_nop;
      rob_13_isComplete <= 1'b0;
      rob_13_branchResult_targetPC <= 32'h00000000;
      rob_13_branchResult_branchResult <= 1'b0;
      rob_13_branchResult_predictFail <= 1'b0;
      rob_13_exceptionInfo_exception <= 1'b0;
      rob_13_exceptionInfo_eCode <= 6'h00;
      rob_13_exceptionInfo_eSubCode <= 1'b0;
      rob_13_valid <= 1'b0;
      rob_14_pc <= 32'h00000000;
      rob_14_ard <= 5'h00;
      rob_14_prd <= 6'h00;
      rob_14_pprd <= 6'h00;
      rob_14_specialOp <= ROBSpecialOp_nop;
      rob_14_isComplete <= 1'b0;
      rob_14_branchResult_targetPC <= 32'h00000000;
      rob_14_branchResult_branchResult <= 1'b0;
      rob_14_branchResult_predictFail <= 1'b0;
      rob_14_exceptionInfo_exception <= 1'b0;
      rob_14_exceptionInfo_eCode <= 6'h00;
      rob_14_exceptionInfo_eSubCode <= 1'b0;
      rob_14_valid <= 1'b0;
      rob_15_pc <= 32'h00000000;
      rob_15_ard <= 5'h00;
      rob_15_prd <= 6'h00;
      rob_15_pprd <= 6'h00;
      rob_15_specialOp <= ROBSpecialOp_nop;
      rob_15_isComplete <= 1'b0;
      rob_15_branchResult_targetPC <= 32'h00000000;
      rob_15_branchResult_branchResult <= 1'b0;
      rob_15_branchResult_predictFail <= 1'b0;
      rob_15_exceptionInfo_exception <= 1'b0;
      rob_15_exceptionInfo_eCode <= 6'h00;
      rob_15_exceptionInfo_eSubCode <= 1'b0;
      rob_15_valid <= 1'b0;
      rob_16_pc <= 32'h00000000;
      rob_16_ard <= 5'h00;
      rob_16_prd <= 6'h00;
      rob_16_pprd <= 6'h00;
      rob_16_specialOp <= ROBSpecialOp_nop;
      rob_16_isComplete <= 1'b0;
      rob_16_branchResult_targetPC <= 32'h00000000;
      rob_16_branchResult_branchResult <= 1'b0;
      rob_16_branchResult_predictFail <= 1'b0;
      rob_16_exceptionInfo_exception <= 1'b0;
      rob_16_exceptionInfo_eCode <= 6'h00;
      rob_16_exceptionInfo_eSubCode <= 1'b0;
      rob_16_valid <= 1'b0;
      rob_17_pc <= 32'h00000000;
      rob_17_ard <= 5'h00;
      rob_17_prd <= 6'h00;
      rob_17_pprd <= 6'h00;
      rob_17_specialOp <= ROBSpecialOp_nop;
      rob_17_isComplete <= 1'b0;
      rob_17_branchResult_targetPC <= 32'h00000000;
      rob_17_branchResult_branchResult <= 1'b0;
      rob_17_branchResult_predictFail <= 1'b0;
      rob_17_exceptionInfo_exception <= 1'b0;
      rob_17_exceptionInfo_eCode <= 6'h00;
      rob_17_exceptionInfo_eSubCode <= 1'b0;
      rob_17_valid <= 1'b0;
      rob_18_pc <= 32'h00000000;
      rob_18_ard <= 5'h00;
      rob_18_prd <= 6'h00;
      rob_18_pprd <= 6'h00;
      rob_18_specialOp <= ROBSpecialOp_nop;
      rob_18_isComplete <= 1'b0;
      rob_18_branchResult_targetPC <= 32'h00000000;
      rob_18_branchResult_branchResult <= 1'b0;
      rob_18_branchResult_predictFail <= 1'b0;
      rob_18_exceptionInfo_exception <= 1'b0;
      rob_18_exceptionInfo_eCode <= 6'h00;
      rob_18_exceptionInfo_eSubCode <= 1'b0;
      rob_18_valid <= 1'b0;
      rob_19_pc <= 32'h00000000;
      rob_19_ard <= 5'h00;
      rob_19_prd <= 6'h00;
      rob_19_pprd <= 6'h00;
      rob_19_specialOp <= ROBSpecialOp_nop;
      rob_19_isComplete <= 1'b0;
      rob_19_branchResult_targetPC <= 32'h00000000;
      rob_19_branchResult_branchResult <= 1'b0;
      rob_19_branchResult_predictFail <= 1'b0;
      rob_19_exceptionInfo_exception <= 1'b0;
      rob_19_exceptionInfo_eCode <= 6'h00;
      rob_19_exceptionInfo_eSubCode <= 1'b0;
      rob_19_valid <= 1'b0;
      rob_20_pc <= 32'h00000000;
      rob_20_ard <= 5'h00;
      rob_20_prd <= 6'h00;
      rob_20_pprd <= 6'h00;
      rob_20_specialOp <= ROBSpecialOp_nop;
      rob_20_isComplete <= 1'b0;
      rob_20_branchResult_targetPC <= 32'h00000000;
      rob_20_branchResult_branchResult <= 1'b0;
      rob_20_branchResult_predictFail <= 1'b0;
      rob_20_exceptionInfo_exception <= 1'b0;
      rob_20_exceptionInfo_eCode <= 6'h00;
      rob_20_exceptionInfo_eSubCode <= 1'b0;
      rob_20_valid <= 1'b0;
      rob_21_pc <= 32'h00000000;
      rob_21_ard <= 5'h00;
      rob_21_prd <= 6'h00;
      rob_21_pprd <= 6'h00;
      rob_21_specialOp <= ROBSpecialOp_nop;
      rob_21_isComplete <= 1'b0;
      rob_21_branchResult_targetPC <= 32'h00000000;
      rob_21_branchResult_branchResult <= 1'b0;
      rob_21_branchResult_predictFail <= 1'b0;
      rob_21_exceptionInfo_exception <= 1'b0;
      rob_21_exceptionInfo_eCode <= 6'h00;
      rob_21_exceptionInfo_eSubCode <= 1'b0;
      rob_21_valid <= 1'b0;
      rob_22_pc <= 32'h00000000;
      rob_22_ard <= 5'h00;
      rob_22_prd <= 6'h00;
      rob_22_pprd <= 6'h00;
      rob_22_specialOp <= ROBSpecialOp_nop;
      rob_22_isComplete <= 1'b0;
      rob_22_branchResult_targetPC <= 32'h00000000;
      rob_22_branchResult_branchResult <= 1'b0;
      rob_22_branchResult_predictFail <= 1'b0;
      rob_22_exceptionInfo_exception <= 1'b0;
      rob_22_exceptionInfo_eCode <= 6'h00;
      rob_22_exceptionInfo_eSubCode <= 1'b0;
      rob_22_valid <= 1'b0;
      rob_23_pc <= 32'h00000000;
      rob_23_ard <= 5'h00;
      rob_23_prd <= 6'h00;
      rob_23_pprd <= 6'h00;
      rob_23_specialOp <= ROBSpecialOp_nop;
      rob_23_isComplete <= 1'b0;
      rob_23_branchResult_targetPC <= 32'h00000000;
      rob_23_branchResult_branchResult <= 1'b0;
      rob_23_branchResult_predictFail <= 1'b0;
      rob_23_exceptionInfo_exception <= 1'b0;
      rob_23_exceptionInfo_eCode <= 6'h00;
      rob_23_exceptionInfo_eSubCode <= 1'b0;
      rob_23_valid <= 1'b0;
      rob_24_pc <= 32'h00000000;
      rob_24_ard <= 5'h00;
      rob_24_prd <= 6'h00;
      rob_24_pprd <= 6'h00;
      rob_24_specialOp <= ROBSpecialOp_nop;
      rob_24_isComplete <= 1'b0;
      rob_24_branchResult_targetPC <= 32'h00000000;
      rob_24_branchResult_branchResult <= 1'b0;
      rob_24_branchResult_predictFail <= 1'b0;
      rob_24_exceptionInfo_exception <= 1'b0;
      rob_24_exceptionInfo_eCode <= 6'h00;
      rob_24_exceptionInfo_eSubCode <= 1'b0;
      rob_24_valid <= 1'b0;
      rob_25_pc <= 32'h00000000;
      rob_25_ard <= 5'h00;
      rob_25_prd <= 6'h00;
      rob_25_pprd <= 6'h00;
      rob_25_specialOp <= ROBSpecialOp_nop;
      rob_25_isComplete <= 1'b0;
      rob_25_branchResult_targetPC <= 32'h00000000;
      rob_25_branchResult_branchResult <= 1'b0;
      rob_25_branchResult_predictFail <= 1'b0;
      rob_25_exceptionInfo_exception <= 1'b0;
      rob_25_exceptionInfo_eCode <= 6'h00;
      rob_25_exceptionInfo_eSubCode <= 1'b0;
      rob_25_valid <= 1'b0;
      rob_26_pc <= 32'h00000000;
      rob_26_ard <= 5'h00;
      rob_26_prd <= 6'h00;
      rob_26_pprd <= 6'h00;
      rob_26_specialOp <= ROBSpecialOp_nop;
      rob_26_isComplete <= 1'b0;
      rob_26_branchResult_targetPC <= 32'h00000000;
      rob_26_branchResult_branchResult <= 1'b0;
      rob_26_branchResult_predictFail <= 1'b0;
      rob_26_exceptionInfo_exception <= 1'b0;
      rob_26_exceptionInfo_eCode <= 6'h00;
      rob_26_exceptionInfo_eSubCode <= 1'b0;
      rob_26_valid <= 1'b0;
      rob_27_pc <= 32'h00000000;
      rob_27_ard <= 5'h00;
      rob_27_prd <= 6'h00;
      rob_27_pprd <= 6'h00;
      rob_27_specialOp <= ROBSpecialOp_nop;
      rob_27_isComplete <= 1'b0;
      rob_27_branchResult_targetPC <= 32'h00000000;
      rob_27_branchResult_branchResult <= 1'b0;
      rob_27_branchResult_predictFail <= 1'b0;
      rob_27_exceptionInfo_exception <= 1'b0;
      rob_27_exceptionInfo_eCode <= 6'h00;
      rob_27_exceptionInfo_eSubCode <= 1'b0;
      rob_27_valid <= 1'b0;
      rob_28_pc <= 32'h00000000;
      rob_28_ard <= 5'h00;
      rob_28_prd <= 6'h00;
      rob_28_pprd <= 6'h00;
      rob_28_specialOp <= ROBSpecialOp_nop;
      rob_28_isComplete <= 1'b0;
      rob_28_branchResult_targetPC <= 32'h00000000;
      rob_28_branchResult_branchResult <= 1'b0;
      rob_28_branchResult_predictFail <= 1'b0;
      rob_28_exceptionInfo_exception <= 1'b0;
      rob_28_exceptionInfo_eCode <= 6'h00;
      rob_28_exceptionInfo_eSubCode <= 1'b0;
      rob_28_valid <= 1'b0;
      rob_29_pc <= 32'h00000000;
      rob_29_ard <= 5'h00;
      rob_29_prd <= 6'h00;
      rob_29_pprd <= 6'h00;
      rob_29_specialOp <= ROBSpecialOp_nop;
      rob_29_isComplete <= 1'b0;
      rob_29_branchResult_targetPC <= 32'h00000000;
      rob_29_branchResult_branchResult <= 1'b0;
      rob_29_branchResult_predictFail <= 1'b0;
      rob_29_exceptionInfo_exception <= 1'b0;
      rob_29_exceptionInfo_eCode <= 6'h00;
      rob_29_exceptionInfo_eSubCode <= 1'b0;
      rob_29_valid <= 1'b0;
      rob_30_pc <= 32'h00000000;
      rob_30_ard <= 5'h00;
      rob_30_prd <= 6'h00;
      rob_30_pprd <= 6'h00;
      rob_30_specialOp <= ROBSpecialOp_nop;
      rob_30_isComplete <= 1'b0;
      rob_30_branchResult_targetPC <= 32'h00000000;
      rob_30_branchResult_branchResult <= 1'b0;
      rob_30_branchResult_predictFail <= 1'b0;
      rob_30_exceptionInfo_exception <= 1'b0;
      rob_30_exceptionInfo_eCode <= 6'h00;
      rob_30_exceptionInfo_eSubCode <= 1'b0;
      rob_30_valid <= 1'b0;
      rob_31_pc <= 32'h00000000;
      rob_31_ard <= 5'h00;
      rob_31_prd <= 6'h00;
      rob_31_pprd <= 6'h00;
      rob_31_specialOp <= ROBSpecialOp_nop;
      rob_31_isComplete <= 1'b0;
      rob_31_branchResult_targetPC <= 32'h00000000;
      rob_31_branchResult_branchResult <= 1'b0;
      rob_31_branchResult_predictFail <= 1'b0;
      rob_31_exceptionInfo_exception <= 1'b0;
      rob_31_exceptionInfo_eCode <= 6'h00;
      rob_31_exceptionInfo_eSubCode <= 1'b0;
      rob_31_valid <= 1'b0;
      head_0 <= 5'h00;
      head_1 <= 5'h01;
      tail_0 <= 5'h00;
      tail_1 <= 5'h01;
      delayedFlush <= 1'b0;
      stageReg_availROBMask <= 2'b00;
      stageReg_retireARAT_0_ard <= 5'h00;
      stageReg_retireARAT_0_prd <= 6'h00;
      stageReg_retireARAT_0_wen <= 1'b0;
      stageReg_retireARAT_1_ard <= 5'h00;
      stageReg_retireARAT_1_prd <= 6'h00;
      stageReg_retireARAT_1_wen <= 1'b0;
      stageReg_freePRFIdx_0 <= 6'h00;
      stageReg_freePRFIdx_1 <= 6'h00;
      stageReg_freePRFNum <= 2'b00;
      stageReg_retireROBIdx_0 <= 5'h00;
      stageReg_retireROBIdx_1 <= 5'h00;
      stageReg_retireEn_0 <= 1'b0;
      stageReg_retireEn_1 <= 1'b0;
      stageReg_wakeupMem <= 1'b0;
      stageReg_retireLLBitUpdate <= 1'b0;
      stageReg_retireWriteCSR <= 1'b0;
      stageReg_retireERTN <= 1'b0;
      stageReg_retireNormalException <= 1'b0;
      stageReg_retireTLBRException <= 1'b0;
      stageReg_retireEPC <= 32'h00000000;
      stageReg_retireEROBIdx <= 5'h00;
      stageReg_retireECode <= 6'h00;
      stageReg_retireESubCode <= 1'b0;
      stageReg_updateBPU_0_pc <= 32'h00000000;
      stageReg_updateBPU_0_isJumpInst <= 1'b0;
      stageReg_updateBPU_0_taken <= 1'b0;
      stageReg_updateBPU_0_predictFail <= 1'b0;
      stageReg_updateBPU_0_target <= 32'h00000000;
      stageReg_updateBPU_1_pc <= 32'h00000000;
      stageReg_updateBPU_1_isJumpInst <= 1'b0;
      stageReg_updateBPU_1_taken <= 1'b0;
      stageReg_updateBPU_1_predictFail <= 1'b0;
      stageReg_updateBPU_1_target <= 32'h00000000;
      stageReg_flush <= 1'b0;
      stageReg_redirectPC <= 32'h00000000;
    end else begin
      rob_0_valid <= (((|_zz_rob_0_isComplete_1) || io_flush) ? 1'b0 : (rob_0_valid || (|_zz_rob_0_valid)));
      rob_0_isComplete <= (((|_zz_rob_0_isComplete_1) || io_flush) ? 1'b0 : (rob_0_isComplete || (|_zz_rob_0_isComplete)));
      rob_1_valid <= (((|_zz_rob_1_isComplete_1) || io_flush) ? 1'b0 : (rob_1_valid || (|_zz_rob_1_valid)));
      rob_1_isComplete <= (((|_zz_rob_1_isComplete_1) || io_flush) ? 1'b0 : (rob_1_isComplete || (|_zz_rob_1_isComplete)));
      rob_2_valid <= (((|_zz_rob_2_isComplete_1) || io_flush) ? 1'b0 : (rob_2_valid || (|_zz_rob_2_valid)));
      rob_2_isComplete <= (((|_zz_rob_2_isComplete_1) || io_flush) ? 1'b0 : (rob_2_isComplete || (|_zz_rob_2_isComplete)));
      rob_3_valid <= (((|_zz_rob_3_isComplete_1) || io_flush) ? 1'b0 : (rob_3_valid || (|_zz_rob_3_valid)));
      rob_3_isComplete <= (((|_zz_rob_3_isComplete_1) || io_flush) ? 1'b0 : (rob_3_isComplete || (|_zz_rob_3_isComplete)));
      rob_4_valid <= (((|_zz_rob_4_isComplete_1) || io_flush) ? 1'b0 : (rob_4_valid || (|_zz_rob_4_valid)));
      rob_4_isComplete <= (((|_zz_rob_4_isComplete_1) || io_flush) ? 1'b0 : (rob_4_isComplete || (|_zz_rob_4_isComplete)));
      rob_5_valid <= (((|_zz_rob_5_isComplete_1) || io_flush) ? 1'b0 : (rob_5_valid || (|_zz_rob_5_valid)));
      rob_5_isComplete <= (((|_zz_rob_5_isComplete_1) || io_flush) ? 1'b0 : (rob_5_isComplete || (|_zz_rob_5_isComplete)));
      rob_6_valid <= (((|_zz_rob_6_isComplete_1) || io_flush) ? 1'b0 : (rob_6_valid || (|_zz_rob_6_valid)));
      rob_6_isComplete <= (((|_zz_rob_6_isComplete_1) || io_flush) ? 1'b0 : (rob_6_isComplete || (|_zz_rob_6_isComplete)));
      rob_7_valid <= (((|_zz_rob_7_isComplete_1) || io_flush) ? 1'b0 : (rob_7_valid || (|_zz_rob_7_valid)));
      rob_7_isComplete <= (((|_zz_rob_7_isComplete_1) || io_flush) ? 1'b0 : (rob_7_isComplete || (|_zz_rob_7_isComplete)));
      rob_8_valid <= (((|_zz_rob_8_isComplete_1) || io_flush) ? 1'b0 : (rob_8_valid || (|_zz_rob_8_valid)));
      rob_8_isComplete <= (((|_zz_rob_8_isComplete_1) || io_flush) ? 1'b0 : (rob_8_isComplete || (|_zz_rob_8_isComplete)));
      rob_9_valid <= (((|_zz_rob_9_isComplete_1) || io_flush) ? 1'b0 : (rob_9_valid || (|_zz_rob_9_valid)));
      rob_9_isComplete <= (((|_zz_rob_9_isComplete_1) || io_flush) ? 1'b0 : (rob_9_isComplete || (|_zz_rob_9_isComplete)));
      rob_10_valid <= (((|_zz_rob_10_isComplete_1) || io_flush) ? 1'b0 : (rob_10_valid || (|_zz_rob_10_valid)));
      rob_10_isComplete <= (((|_zz_rob_10_isComplete_1) || io_flush) ? 1'b0 : (rob_10_isComplete || (|_zz_rob_10_isComplete)));
      rob_11_valid <= (((|_zz_rob_11_isComplete_1) || io_flush) ? 1'b0 : (rob_11_valid || (|_zz_rob_11_valid)));
      rob_11_isComplete <= (((|_zz_rob_11_isComplete_1) || io_flush) ? 1'b0 : (rob_11_isComplete || (|_zz_rob_11_isComplete)));
      rob_12_valid <= (((|_zz_rob_12_isComplete_1) || io_flush) ? 1'b0 : (rob_12_valid || (|_zz_rob_12_valid)));
      rob_12_isComplete <= (((|_zz_rob_12_isComplete_1) || io_flush) ? 1'b0 : (rob_12_isComplete || (|_zz_rob_12_isComplete)));
      rob_13_valid <= (((|_zz_rob_13_isComplete_1) || io_flush) ? 1'b0 : (rob_13_valid || (|_zz_rob_13_valid)));
      rob_13_isComplete <= (((|_zz_rob_13_isComplete_1) || io_flush) ? 1'b0 : (rob_13_isComplete || (|_zz_rob_13_isComplete)));
      rob_14_valid <= (((|_zz_rob_14_isComplete_1) || io_flush) ? 1'b0 : (rob_14_valid || (|_zz_rob_14_valid)));
      rob_14_isComplete <= (((|_zz_rob_14_isComplete_1) || io_flush) ? 1'b0 : (rob_14_isComplete || (|_zz_rob_14_isComplete)));
      rob_15_valid <= (((|_zz_rob_15_isComplete_1) || io_flush) ? 1'b0 : (rob_15_valid || (|_zz_rob_15_valid)));
      rob_15_isComplete <= (((|_zz_rob_15_isComplete_1) || io_flush) ? 1'b0 : (rob_15_isComplete || (|_zz_rob_15_isComplete)));
      rob_16_valid <= (((|_zz_rob_16_isComplete_1) || io_flush) ? 1'b0 : (rob_16_valid || (|_zz_rob_16_valid)));
      rob_16_isComplete <= (((|_zz_rob_16_isComplete_1) || io_flush) ? 1'b0 : (rob_16_isComplete || (|_zz_rob_16_isComplete)));
      rob_17_valid <= (((|_zz_rob_17_isComplete_1) || io_flush) ? 1'b0 : (rob_17_valid || (|_zz_rob_17_valid)));
      rob_17_isComplete <= (((|_zz_rob_17_isComplete_1) || io_flush) ? 1'b0 : (rob_17_isComplete || (|_zz_rob_17_isComplete)));
      rob_18_valid <= (((|_zz_rob_18_isComplete_1) || io_flush) ? 1'b0 : (rob_18_valid || (|_zz_rob_18_valid)));
      rob_18_isComplete <= (((|_zz_rob_18_isComplete_1) || io_flush) ? 1'b0 : (rob_18_isComplete || (|_zz_rob_18_isComplete)));
      rob_19_valid <= (((|_zz_rob_19_isComplete_1) || io_flush) ? 1'b0 : (rob_19_valid || (|_zz_rob_19_valid)));
      rob_19_isComplete <= (((|_zz_rob_19_isComplete_1) || io_flush) ? 1'b0 : (rob_19_isComplete || (|_zz_rob_19_isComplete)));
      rob_20_valid <= (((|_zz_rob_20_isComplete_1) || io_flush) ? 1'b0 : (rob_20_valid || (|_zz_rob_20_valid)));
      rob_20_isComplete <= (((|_zz_rob_20_isComplete_1) || io_flush) ? 1'b0 : (rob_20_isComplete || (|_zz_rob_20_isComplete)));
      rob_21_valid <= (((|_zz_rob_21_isComplete_1) || io_flush) ? 1'b0 : (rob_21_valid || (|_zz_rob_21_valid)));
      rob_21_isComplete <= (((|_zz_rob_21_isComplete_1) || io_flush) ? 1'b0 : (rob_21_isComplete || (|_zz_rob_21_isComplete)));
      rob_22_valid <= (((|_zz_rob_22_isComplete_1) || io_flush) ? 1'b0 : (rob_22_valid || (|_zz_rob_22_valid)));
      rob_22_isComplete <= (((|_zz_rob_22_isComplete_1) || io_flush) ? 1'b0 : (rob_22_isComplete || (|_zz_rob_22_isComplete)));
      rob_23_valid <= (((|_zz_rob_23_isComplete_1) || io_flush) ? 1'b0 : (rob_23_valid || (|_zz_rob_23_valid)));
      rob_23_isComplete <= (((|_zz_rob_23_isComplete_1) || io_flush) ? 1'b0 : (rob_23_isComplete || (|_zz_rob_23_isComplete)));
      rob_24_valid <= (((|_zz_rob_24_isComplete_1) || io_flush) ? 1'b0 : (rob_24_valid || (|_zz_rob_24_valid)));
      rob_24_isComplete <= (((|_zz_rob_24_isComplete_1) || io_flush) ? 1'b0 : (rob_24_isComplete || (|_zz_rob_24_isComplete)));
      rob_25_valid <= (((|_zz_rob_25_isComplete_1) || io_flush) ? 1'b0 : (rob_25_valid || (|_zz_rob_25_valid)));
      rob_25_isComplete <= (((|_zz_rob_25_isComplete_1) || io_flush) ? 1'b0 : (rob_25_isComplete || (|_zz_rob_25_isComplete)));
      rob_26_valid <= (((|_zz_rob_26_isComplete_1) || io_flush) ? 1'b0 : (rob_26_valid || (|_zz_rob_26_valid)));
      rob_26_isComplete <= (((|_zz_rob_26_isComplete_1) || io_flush) ? 1'b0 : (rob_26_isComplete || (|_zz_rob_26_isComplete)));
      rob_27_valid <= (((|_zz_rob_27_isComplete_1) || io_flush) ? 1'b0 : (rob_27_valid || (|_zz_rob_27_valid)));
      rob_27_isComplete <= (((|_zz_rob_27_isComplete_1) || io_flush) ? 1'b0 : (rob_27_isComplete || (|_zz_rob_27_isComplete)));
      rob_28_valid <= (((|_zz_rob_28_isComplete_1) || io_flush) ? 1'b0 : (rob_28_valid || (|_zz_rob_28_valid)));
      rob_28_isComplete <= (((|_zz_rob_28_isComplete_1) || io_flush) ? 1'b0 : (rob_28_isComplete || (|_zz_rob_28_isComplete)));
      rob_29_valid <= (((|_zz_rob_29_isComplete_1) || io_flush) ? 1'b0 : (rob_29_valid || (|_zz_rob_29_valid)));
      rob_29_isComplete <= (((|_zz_rob_29_isComplete_1) || io_flush) ? 1'b0 : (rob_29_isComplete || (|_zz_rob_29_isComplete)));
      rob_30_valid <= (((|_zz_rob_30_isComplete_1) || io_flush) ? 1'b0 : (rob_30_valid || (|_zz_rob_30_valid)));
      rob_30_isComplete <= (((|_zz_rob_30_isComplete_1) || io_flush) ? 1'b0 : (rob_30_isComplete || (|_zz_rob_30_isComplete)));
      rob_31_valid <= (((|_zz_rob_31_isComplete_1) || io_flush) ? 1'b0 : (rob_31_valid || (|_zz_rob_31_valid)));
      rob_31_isComplete <= (((|_zz_rob_31_isComplete_1) || io_flush) ? 1'b0 : (rob_31_isComplete || (|_zz_rob_31_isComplete)));
      if(when_ROB_l76) begin
        if(_zz_2) begin
          rob_0_pc <= io_dispatch_pc_0;
        end
        if(_zz_3) begin
          rob_1_pc <= io_dispatch_pc_0;
        end
        if(_zz_4) begin
          rob_2_pc <= io_dispatch_pc_0;
        end
        if(_zz_5) begin
          rob_3_pc <= io_dispatch_pc_0;
        end
        if(_zz_6) begin
          rob_4_pc <= io_dispatch_pc_0;
        end
        if(_zz_7) begin
          rob_5_pc <= io_dispatch_pc_0;
        end
        if(_zz_8) begin
          rob_6_pc <= io_dispatch_pc_0;
        end
        if(_zz_9) begin
          rob_7_pc <= io_dispatch_pc_0;
        end
        if(_zz_10) begin
          rob_8_pc <= io_dispatch_pc_0;
        end
        if(_zz_11) begin
          rob_9_pc <= io_dispatch_pc_0;
        end
        if(_zz_12) begin
          rob_10_pc <= io_dispatch_pc_0;
        end
        if(_zz_13) begin
          rob_11_pc <= io_dispatch_pc_0;
        end
        if(_zz_14) begin
          rob_12_pc <= io_dispatch_pc_0;
        end
        if(_zz_15) begin
          rob_13_pc <= io_dispatch_pc_0;
        end
        if(_zz_16) begin
          rob_14_pc <= io_dispatch_pc_0;
        end
        if(_zz_17) begin
          rob_15_pc <= io_dispatch_pc_0;
        end
        if(_zz_18) begin
          rob_16_pc <= io_dispatch_pc_0;
        end
        if(_zz_19) begin
          rob_17_pc <= io_dispatch_pc_0;
        end
        if(_zz_20) begin
          rob_18_pc <= io_dispatch_pc_0;
        end
        if(_zz_21) begin
          rob_19_pc <= io_dispatch_pc_0;
        end
        if(_zz_22) begin
          rob_20_pc <= io_dispatch_pc_0;
        end
        if(_zz_23) begin
          rob_21_pc <= io_dispatch_pc_0;
        end
        if(_zz_24) begin
          rob_22_pc <= io_dispatch_pc_0;
        end
        if(_zz_25) begin
          rob_23_pc <= io_dispatch_pc_0;
        end
        if(_zz_26) begin
          rob_24_pc <= io_dispatch_pc_0;
        end
        if(_zz_27) begin
          rob_25_pc <= io_dispatch_pc_0;
        end
        if(_zz_28) begin
          rob_26_pc <= io_dispatch_pc_0;
        end
        if(_zz_29) begin
          rob_27_pc <= io_dispatch_pc_0;
        end
        if(_zz_30) begin
          rob_28_pc <= io_dispatch_pc_0;
        end
        if(_zz_31) begin
          rob_29_pc <= io_dispatch_pc_0;
        end
        if(_zz_32) begin
          rob_30_pc <= io_dispatch_pc_0;
        end
        if(_zz_33) begin
          rob_31_pc <= io_dispatch_pc_0;
        end
        if(_zz_2) begin
          rob_0_ard <= io_dispatch_ard_0;
        end
        if(_zz_3) begin
          rob_1_ard <= io_dispatch_ard_0;
        end
        if(_zz_4) begin
          rob_2_ard <= io_dispatch_ard_0;
        end
        if(_zz_5) begin
          rob_3_ard <= io_dispatch_ard_0;
        end
        if(_zz_6) begin
          rob_4_ard <= io_dispatch_ard_0;
        end
        if(_zz_7) begin
          rob_5_ard <= io_dispatch_ard_0;
        end
        if(_zz_8) begin
          rob_6_ard <= io_dispatch_ard_0;
        end
        if(_zz_9) begin
          rob_7_ard <= io_dispatch_ard_0;
        end
        if(_zz_10) begin
          rob_8_ard <= io_dispatch_ard_0;
        end
        if(_zz_11) begin
          rob_9_ard <= io_dispatch_ard_0;
        end
        if(_zz_12) begin
          rob_10_ard <= io_dispatch_ard_0;
        end
        if(_zz_13) begin
          rob_11_ard <= io_dispatch_ard_0;
        end
        if(_zz_14) begin
          rob_12_ard <= io_dispatch_ard_0;
        end
        if(_zz_15) begin
          rob_13_ard <= io_dispatch_ard_0;
        end
        if(_zz_16) begin
          rob_14_ard <= io_dispatch_ard_0;
        end
        if(_zz_17) begin
          rob_15_ard <= io_dispatch_ard_0;
        end
        if(_zz_18) begin
          rob_16_ard <= io_dispatch_ard_0;
        end
        if(_zz_19) begin
          rob_17_ard <= io_dispatch_ard_0;
        end
        if(_zz_20) begin
          rob_18_ard <= io_dispatch_ard_0;
        end
        if(_zz_21) begin
          rob_19_ard <= io_dispatch_ard_0;
        end
        if(_zz_22) begin
          rob_20_ard <= io_dispatch_ard_0;
        end
        if(_zz_23) begin
          rob_21_ard <= io_dispatch_ard_0;
        end
        if(_zz_24) begin
          rob_22_ard <= io_dispatch_ard_0;
        end
        if(_zz_25) begin
          rob_23_ard <= io_dispatch_ard_0;
        end
        if(_zz_26) begin
          rob_24_ard <= io_dispatch_ard_0;
        end
        if(_zz_27) begin
          rob_25_ard <= io_dispatch_ard_0;
        end
        if(_zz_28) begin
          rob_26_ard <= io_dispatch_ard_0;
        end
        if(_zz_29) begin
          rob_27_ard <= io_dispatch_ard_0;
        end
        if(_zz_30) begin
          rob_28_ard <= io_dispatch_ard_0;
        end
        if(_zz_31) begin
          rob_29_ard <= io_dispatch_ard_0;
        end
        if(_zz_32) begin
          rob_30_ard <= io_dispatch_ard_0;
        end
        if(_zz_33) begin
          rob_31_ard <= io_dispatch_ard_0;
        end
        if(_zz_2) begin
          rob_0_prd <= io_dispatch_prd_0;
        end
        if(_zz_3) begin
          rob_1_prd <= io_dispatch_prd_0;
        end
        if(_zz_4) begin
          rob_2_prd <= io_dispatch_prd_0;
        end
        if(_zz_5) begin
          rob_3_prd <= io_dispatch_prd_0;
        end
        if(_zz_6) begin
          rob_4_prd <= io_dispatch_prd_0;
        end
        if(_zz_7) begin
          rob_5_prd <= io_dispatch_prd_0;
        end
        if(_zz_8) begin
          rob_6_prd <= io_dispatch_prd_0;
        end
        if(_zz_9) begin
          rob_7_prd <= io_dispatch_prd_0;
        end
        if(_zz_10) begin
          rob_8_prd <= io_dispatch_prd_0;
        end
        if(_zz_11) begin
          rob_9_prd <= io_dispatch_prd_0;
        end
        if(_zz_12) begin
          rob_10_prd <= io_dispatch_prd_0;
        end
        if(_zz_13) begin
          rob_11_prd <= io_dispatch_prd_0;
        end
        if(_zz_14) begin
          rob_12_prd <= io_dispatch_prd_0;
        end
        if(_zz_15) begin
          rob_13_prd <= io_dispatch_prd_0;
        end
        if(_zz_16) begin
          rob_14_prd <= io_dispatch_prd_0;
        end
        if(_zz_17) begin
          rob_15_prd <= io_dispatch_prd_0;
        end
        if(_zz_18) begin
          rob_16_prd <= io_dispatch_prd_0;
        end
        if(_zz_19) begin
          rob_17_prd <= io_dispatch_prd_0;
        end
        if(_zz_20) begin
          rob_18_prd <= io_dispatch_prd_0;
        end
        if(_zz_21) begin
          rob_19_prd <= io_dispatch_prd_0;
        end
        if(_zz_22) begin
          rob_20_prd <= io_dispatch_prd_0;
        end
        if(_zz_23) begin
          rob_21_prd <= io_dispatch_prd_0;
        end
        if(_zz_24) begin
          rob_22_prd <= io_dispatch_prd_0;
        end
        if(_zz_25) begin
          rob_23_prd <= io_dispatch_prd_0;
        end
        if(_zz_26) begin
          rob_24_prd <= io_dispatch_prd_0;
        end
        if(_zz_27) begin
          rob_25_prd <= io_dispatch_prd_0;
        end
        if(_zz_28) begin
          rob_26_prd <= io_dispatch_prd_0;
        end
        if(_zz_29) begin
          rob_27_prd <= io_dispatch_prd_0;
        end
        if(_zz_30) begin
          rob_28_prd <= io_dispatch_prd_0;
        end
        if(_zz_31) begin
          rob_29_prd <= io_dispatch_prd_0;
        end
        if(_zz_32) begin
          rob_30_prd <= io_dispatch_prd_0;
        end
        if(_zz_33) begin
          rob_31_prd <= io_dispatch_prd_0;
        end
        if(_zz_2) begin
          rob_0_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_3) begin
          rob_1_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_4) begin
          rob_2_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_5) begin
          rob_3_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_6) begin
          rob_4_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_7) begin
          rob_5_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_8) begin
          rob_6_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_9) begin
          rob_7_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_10) begin
          rob_8_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_11) begin
          rob_9_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_12) begin
          rob_10_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_13) begin
          rob_11_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_14) begin
          rob_12_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_15) begin
          rob_13_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_16) begin
          rob_14_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_17) begin
          rob_15_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_18) begin
          rob_16_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_19) begin
          rob_17_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_20) begin
          rob_18_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_21) begin
          rob_19_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_22) begin
          rob_20_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_23) begin
          rob_21_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_24) begin
          rob_22_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_25) begin
          rob_23_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_26) begin
          rob_24_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_27) begin
          rob_25_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_28) begin
          rob_26_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_29) begin
          rob_27_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_30) begin
          rob_28_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_31) begin
          rob_29_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_32) begin
          rob_30_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_33) begin
          rob_31_pprd <= io_dispatch_pprd_0;
        end
        if(_zz_2) begin
          rob_0_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_3) begin
          rob_1_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_4) begin
          rob_2_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_5) begin
          rob_3_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_6) begin
          rob_4_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_7) begin
          rob_5_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_8) begin
          rob_6_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_9) begin
          rob_7_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_10) begin
          rob_8_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_11) begin
          rob_9_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_12) begin
          rob_10_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_13) begin
          rob_11_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_14) begin
          rob_12_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_15) begin
          rob_13_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_16) begin
          rob_14_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_17) begin
          rob_15_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_18) begin
          rob_16_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_19) begin
          rob_17_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_20) begin
          rob_18_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_21) begin
          rob_19_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_22) begin
          rob_20_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_23) begin
          rob_21_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_24) begin
          rob_22_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_25) begin
          rob_23_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_26) begin
          rob_24_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_27) begin
          rob_25_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_28) begin
          rob_26_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_29) begin
          rob_27_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_30) begin
          rob_28_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_31) begin
          rob_29_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_32) begin
          rob_30_specialOp <= io_dispatch_specialOp_0;
        end
        if(_zz_33) begin
          rob_31_specialOp <= io_dispatch_specialOp_0;
        end
      end
      tail_0 <= (io_flush ? 5'h00 : _zz_tail_0);
      if(when_ROB_l76_1) begin
        if(_zz_35) begin
          rob_0_pc <= io_dispatch_pc_1;
        end
        if(_zz_36) begin
          rob_1_pc <= io_dispatch_pc_1;
        end
        if(_zz_37) begin
          rob_2_pc <= io_dispatch_pc_1;
        end
        if(_zz_38) begin
          rob_3_pc <= io_dispatch_pc_1;
        end
        if(_zz_39) begin
          rob_4_pc <= io_dispatch_pc_1;
        end
        if(_zz_40) begin
          rob_5_pc <= io_dispatch_pc_1;
        end
        if(_zz_41) begin
          rob_6_pc <= io_dispatch_pc_1;
        end
        if(_zz_42) begin
          rob_7_pc <= io_dispatch_pc_1;
        end
        if(_zz_43) begin
          rob_8_pc <= io_dispatch_pc_1;
        end
        if(_zz_44) begin
          rob_9_pc <= io_dispatch_pc_1;
        end
        if(_zz_45) begin
          rob_10_pc <= io_dispatch_pc_1;
        end
        if(_zz_46) begin
          rob_11_pc <= io_dispatch_pc_1;
        end
        if(_zz_47) begin
          rob_12_pc <= io_dispatch_pc_1;
        end
        if(_zz_48) begin
          rob_13_pc <= io_dispatch_pc_1;
        end
        if(_zz_49) begin
          rob_14_pc <= io_dispatch_pc_1;
        end
        if(_zz_50) begin
          rob_15_pc <= io_dispatch_pc_1;
        end
        if(_zz_51) begin
          rob_16_pc <= io_dispatch_pc_1;
        end
        if(_zz_52) begin
          rob_17_pc <= io_dispatch_pc_1;
        end
        if(_zz_53) begin
          rob_18_pc <= io_dispatch_pc_1;
        end
        if(_zz_54) begin
          rob_19_pc <= io_dispatch_pc_1;
        end
        if(_zz_55) begin
          rob_20_pc <= io_dispatch_pc_1;
        end
        if(_zz_56) begin
          rob_21_pc <= io_dispatch_pc_1;
        end
        if(_zz_57) begin
          rob_22_pc <= io_dispatch_pc_1;
        end
        if(_zz_58) begin
          rob_23_pc <= io_dispatch_pc_1;
        end
        if(_zz_59) begin
          rob_24_pc <= io_dispatch_pc_1;
        end
        if(_zz_60) begin
          rob_25_pc <= io_dispatch_pc_1;
        end
        if(_zz_61) begin
          rob_26_pc <= io_dispatch_pc_1;
        end
        if(_zz_62) begin
          rob_27_pc <= io_dispatch_pc_1;
        end
        if(_zz_63) begin
          rob_28_pc <= io_dispatch_pc_1;
        end
        if(_zz_64) begin
          rob_29_pc <= io_dispatch_pc_1;
        end
        if(_zz_65) begin
          rob_30_pc <= io_dispatch_pc_1;
        end
        if(_zz_66) begin
          rob_31_pc <= io_dispatch_pc_1;
        end
        if(_zz_35) begin
          rob_0_ard <= io_dispatch_ard_1;
        end
        if(_zz_36) begin
          rob_1_ard <= io_dispatch_ard_1;
        end
        if(_zz_37) begin
          rob_2_ard <= io_dispatch_ard_1;
        end
        if(_zz_38) begin
          rob_3_ard <= io_dispatch_ard_1;
        end
        if(_zz_39) begin
          rob_4_ard <= io_dispatch_ard_1;
        end
        if(_zz_40) begin
          rob_5_ard <= io_dispatch_ard_1;
        end
        if(_zz_41) begin
          rob_6_ard <= io_dispatch_ard_1;
        end
        if(_zz_42) begin
          rob_7_ard <= io_dispatch_ard_1;
        end
        if(_zz_43) begin
          rob_8_ard <= io_dispatch_ard_1;
        end
        if(_zz_44) begin
          rob_9_ard <= io_dispatch_ard_1;
        end
        if(_zz_45) begin
          rob_10_ard <= io_dispatch_ard_1;
        end
        if(_zz_46) begin
          rob_11_ard <= io_dispatch_ard_1;
        end
        if(_zz_47) begin
          rob_12_ard <= io_dispatch_ard_1;
        end
        if(_zz_48) begin
          rob_13_ard <= io_dispatch_ard_1;
        end
        if(_zz_49) begin
          rob_14_ard <= io_dispatch_ard_1;
        end
        if(_zz_50) begin
          rob_15_ard <= io_dispatch_ard_1;
        end
        if(_zz_51) begin
          rob_16_ard <= io_dispatch_ard_1;
        end
        if(_zz_52) begin
          rob_17_ard <= io_dispatch_ard_1;
        end
        if(_zz_53) begin
          rob_18_ard <= io_dispatch_ard_1;
        end
        if(_zz_54) begin
          rob_19_ard <= io_dispatch_ard_1;
        end
        if(_zz_55) begin
          rob_20_ard <= io_dispatch_ard_1;
        end
        if(_zz_56) begin
          rob_21_ard <= io_dispatch_ard_1;
        end
        if(_zz_57) begin
          rob_22_ard <= io_dispatch_ard_1;
        end
        if(_zz_58) begin
          rob_23_ard <= io_dispatch_ard_1;
        end
        if(_zz_59) begin
          rob_24_ard <= io_dispatch_ard_1;
        end
        if(_zz_60) begin
          rob_25_ard <= io_dispatch_ard_1;
        end
        if(_zz_61) begin
          rob_26_ard <= io_dispatch_ard_1;
        end
        if(_zz_62) begin
          rob_27_ard <= io_dispatch_ard_1;
        end
        if(_zz_63) begin
          rob_28_ard <= io_dispatch_ard_1;
        end
        if(_zz_64) begin
          rob_29_ard <= io_dispatch_ard_1;
        end
        if(_zz_65) begin
          rob_30_ard <= io_dispatch_ard_1;
        end
        if(_zz_66) begin
          rob_31_ard <= io_dispatch_ard_1;
        end
        if(_zz_35) begin
          rob_0_prd <= io_dispatch_prd_1;
        end
        if(_zz_36) begin
          rob_1_prd <= io_dispatch_prd_1;
        end
        if(_zz_37) begin
          rob_2_prd <= io_dispatch_prd_1;
        end
        if(_zz_38) begin
          rob_3_prd <= io_dispatch_prd_1;
        end
        if(_zz_39) begin
          rob_4_prd <= io_dispatch_prd_1;
        end
        if(_zz_40) begin
          rob_5_prd <= io_dispatch_prd_1;
        end
        if(_zz_41) begin
          rob_6_prd <= io_dispatch_prd_1;
        end
        if(_zz_42) begin
          rob_7_prd <= io_dispatch_prd_1;
        end
        if(_zz_43) begin
          rob_8_prd <= io_dispatch_prd_1;
        end
        if(_zz_44) begin
          rob_9_prd <= io_dispatch_prd_1;
        end
        if(_zz_45) begin
          rob_10_prd <= io_dispatch_prd_1;
        end
        if(_zz_46) begin
          rob_11_prd <= io_dispatch_prd_1;
        end
        if(_zz_47) begin
          rob_12_prd <= io_dispatch_prd_1;
        end
        if(_zz_48) begin
          rob_13_prd <= io_dispatch_prd_1;
        end
        if(_zz_49) begin
          rob_14_prd <= io_dispatch_prd_1;
        end
        if(_zz_50) begin
          rob_15_prd <= io_dispatch_prd_1;
        end
        if(_zz_51) begin
          rob_16_prd <= io_dispatch_prd_1;
        end
        if(_zz_52) begin
          rob_17_prd <= io_dispatch_prd_1;
        end
        if(_zz_53) begin
          rob_18_prd <= io_dispatch_prd_1;
        end
        if(_zz_54) begin
          rob_19_prd <= io_dispatch_prd_1;
        end
        if(_zz_55) begin
          rob_20_prd <= io_dispatch_prd_1;
        end
        if(_zz_56) begin
          rob_21_prd <= io_dispatch_prd_1;
        end
        if(_zz_57) begin
          rob_22_prd <= io_dispatch_prd_1;
        end
        if(_zz_58) begin
          rob_23_prd <= io_dispatch_prd_1;
        end
        if(_zz_59) begin
          rob_24_prd <= io_dispatch_prd_1;
        end
        if(_zz_60) begin
          rob_25_prd <= io_dispatch_prd_1;
        end
        if(_zz_61) begin
          rob_26_prd <= io_dispatch_prd_1;
        end
        if(_zz_62) begin
          rob_27_prd <= io_dispatch_prd_1;
        end
        if(_zz_63) begin
          rob_28_prd <= io_dispatch_prd_1;
        end
        if(_zz_64) begin
          rob_29_prd <= io_dispatch_prd_1;
        end
        if(_zz_65) begin
          rob_30_prd <= io_dispatch_prd_1;
        end
        if(_zz_66) begin
          rob_31_prd <= io_dispatch_prd_1;
        end
        if(_zz_35) begin
          rob_0_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_36) begin
          rob_1_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_37) begin
          rob_2_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_38) begin
          rob_3_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_39) begin
          rob_4_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_40) begin
          rob_5_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_41) begin
          rob_6_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_42) begin
          rob_7_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_43) begin
          rob_8_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_44) begin
          rob_9_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_45) begin
          rob_10_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_46) begin
          rob_11_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_47) begin
          rob_12_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_48) begin
          rob_13_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_49) begin
          rob_14_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_50) begin
          rob_15_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_51) begin
          rob_16_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_52) begin
          rob_17_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_53) begin
          rob_18_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_54) begin
          rob_19_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_55) begin
          rob_20_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_56) begin
          rob_21_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_57) begin
          rob_22_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_58) begin
          rob_23_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_59) begin
          rob_24_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_60) begin
          rob_25_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_61) begin
          rob_26_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_62) begin
          rob_27_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_63) begin
          rob_28_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_64) begin
          rob_29_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_65) begin
          rob_30_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_66) begin
          rob_31_pprd <= io_dispatch_pprd_1;
        end
        if(_zz_35) begin
          rob_0_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_36) begin
          rob_1_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_37) begin
          rob_2_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_38) begin
          rob_3_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_39) begin
          rob_4_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_40) begin
          rob_5_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_41) begin
          rob_6_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_42) begin
          rob_7_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_43) begin
          rob_8_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_44) begin
          rob_9_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_45) begin
          rob_10_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_46) begin
          rob_11_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_47) begin
          rob_12_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_48) begin
          rob_13_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_49) begin
          rob_14_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_50) begin
          rob_15_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_51) begin
          rob_16_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_52) begin
          rob_17_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_53) begin
          rob_18_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_54) begin
          rob_19_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_55) begin
          rob_20_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_56) begin
          rob_21_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_57) begin
          rob_22_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_58) begin
          rob_23_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_59) begin
          rob_24_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_60) begin
          rob_25_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_61) begin
          rob_26_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_62) begin
          rob_27_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_63) begin
          rob_28_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_64) begin
          rob_29_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_65) begin
          rob_30_specialOp <= io_dispatch_specialOp_1;
        end
        if(_zz_66) begin
          rob_31_specialOp <= io_dispatch_specialOp_1;
        end
      end
      tail_1 <= (io_flush ? _zz_tail_1 : _zz_tail_1_2);
      if(io_commit_0_valid) begin
        if(_zz_68) begin
          rob_0_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_69) begin
          rob_1_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_70) begin
          rob_2_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_71) begin
          rob_3_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_72) begin
          rob_4_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_73) begin
          rob_5_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_74) begin
          rob_6_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_75) begin
          rob_7_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_76) begin
          rob_8_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_77) begin
          rob_9_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_78) begin
          rob_10_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_79) begin
          rob_11_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_80) begin
          rob_12_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_81) begin
          rob_13_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_82) begin
          rob_14_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_83) begin
          rob_15_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_84) begin
          rob_16_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_85) begin
          rob_17_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_86) begin
          rob_18_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_87) begin
          rob_19_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_88) begin
          rob_20_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_89) begin
          rob_21_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_90) begin
          rob_22_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_91) begin
          rob_23_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_92) begin
          rob_24_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_93) begin
          rob_25_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_94) begin
          rob_26_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_95) begin
          rob_27_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_96) begin
          rob_28_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_97) begin
          rob_29_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_98) begin
          rob_30_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_99) begin
          rob_31_branchResult_targetPC <= io_commit_0_branchResult_targetPC;
        end
        if(_zz_68) begin
          rob_0_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_69) begin
          rob_1_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_70) begin
          rob_2_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_71) begin
          rob_3_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_72) begin
          rob_4_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_73) begin
          rob_5_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_74) begin
          rob_6_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_75) begin
          rob_7_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_76) begin
          rob_8_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_77) begin
          rob_9_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_78) begin
          rob_10_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_79) begin
          rob_11_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_80) begin
          rob_12_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_81) begin
          rob_13_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_82) begin
          rob_14_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_83) begin
          rob_15_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_84) begin
          rob_16_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_85) begin
          rob_17_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_86) begin
          rob_18_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_87) begin
          rob_19_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_88) begin
          rob_20_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_89) begin
          rob_21_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_90) begin
          rob_22_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_91) begin
          rob_23_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_92) begin
          rob_24_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_93) begin
          rob_25_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_94) begin
          rob_26_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_95) begin
          rob_27_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_96) begin
          rob_28_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_97) begin
          rob_29_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_98) begin
          rob_30_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_99) begin
          rob_31_branchResult_branchResult <= io_commit_0_branchResult_branchResult;
        end
        if(_zz_68) begin
          rob_0_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_69) begin
          rob_1_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_70) begin
          rob_2_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_71) begin
          rob_3_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_72) begin
          rob_4_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_73) begin
          rob_5_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_74) begin
          rob_6_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_75) begin
          rob_7_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_76) begin
          rob_8_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_77) begin
          rob_9_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_78) begin
          rob_10_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_79) begin
          rob_11_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_80) begin
          rob_12_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_81) begin
          rob_13_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_82) begin
          rob_14_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_83) begin
          rob_15_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_84) begin
          rob_16_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_85) begin
          rob_17_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_86) begin
          rob_18_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_87) begin
          rob_19_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_88) begin
          rob_20_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_89) begin
          rob_21_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_90) begin
          rob_22_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_91) begin
          rob_23_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_92) begin
          rob_24_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_93) begin
          rob_25_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_94) begin
          rob_26_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_95) begin
          rob_27_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_96) begin
          rob_28_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_97) begin
          rob_29_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_98) begin
          rob_30_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_99) begin
          rob_31_branchResult_predictFail <= io_commit_0_branchResult_predictFail;
        end
        if(_zz_101) begin
          rob_0_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_102) begin
          rob_1_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_103) begin
          rob_2_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_104) begin
          rob_3_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_105) begin
          rob_4_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_106) begin
          rob_5_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_107) begin
          rob_6_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_108) begin
          rob_7_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_109) begin
          rob_8_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_110) begin
          rob_9_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_111) begin
          rob_10_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_112) begin
          rob_11_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_113) begin
          rob_12_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_114) begin
          rob_13_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_115) begin
          rob_14_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_116) begin
          rob_15_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_117) begin
          rob_16_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_118) begin
          rob_17_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_119) begin
          rob_18_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_120) begin
          rob_19_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_121) begin
          rob_20_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_122) begin
          rob_21_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_123) begin
          rob_22_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_124) begin
          rob_23_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_125) begin
          rob_24_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_126) begin
          rob_25_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_127) begin
          rob_26_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_128) begin
          rob_27_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_129) begin
          rob_28_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_130) begin
          rob_29_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_131) begin
          rob_30_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_132) begin
          rob_31_exceptionInfo_exception <= io_commit_0_exceptionInfo_exception;
        end
        if(_zz_101) begin
          rob_0_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_102) begin
          rob_1_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_103) begin
          rob_2_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_104) begin
          rob_3_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_105) begin
          rob_4_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_106) begin
          rob_5_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_107) begin
          rob_6_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_108) begin
          rob_7_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_109) begin
          rob_8_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_110) begin
          rob_9_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_111) begin
          rob_10_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_112) begin
          rob_11_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_113) begin
          rob_12_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_114) begin
          rob_13_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_115) begin
          rob_14_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_116) begin
          rob_15_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_117) begin
          rob_16_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_118) begin
          rob_17_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_119) begin
          rob_18_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_120) begin
          rob_19_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_121) begin
          rob_20_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_122) begin
          rob_21_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_123) begin
          rob_22_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_124) begin
          rob_23_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_125) begin
          rob_24_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_126) begin
          rob_25_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_127) begin
          rob_26_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_128) begin
          rob_27_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_129) begin
          rob_28_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_130) begin
          rob_29_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_131) begin
          rob_30_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_132) begin
          rob_31_exceptionInfo_eCode <= io_commit_0_exceptionInfo_eCode;
        end
        if(_zz_101) begin
          rob_0_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_102) begin
          rob_1_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_103) begin
          rob_2_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_104) begin
          rob_3_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_105) begin
          rob_4_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_106) begin
          rob_5_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_107) begin
          rob_6_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_108) begin
          rob_7_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_109) begin
          rob_8_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_110) begin
          rob_9_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_111) begin
          rob_10_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_112) begin
          rob_11_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_113) begin
          rob_12_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_114) begin
          rob_13_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_115) begin
          rob_14_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_116) begin
          rob_15_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_117) begin
          rob_16_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_118) begin
          rob_17_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_119) begin
          rob_18_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_120) begin
          rob_19_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_121) begin
          rob_20_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_122) begin
          rob_21_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_123) begin
          rob_22_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_124) begin
          rob_23_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_125) begin
          rob_24_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_126) begin
          rob_25_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_127) begin
          rob_26_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_128) begin
          rob_27_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_129) begin
          rob_28_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_130) begin
          rob_29_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_131) begin
          rob_30_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
        if(_zz_132) begin
          rob_31_exceptionInfo_eSubCode <= io_commit_0_exceptionInfo_eSubCode;
        end
      end
      if(io_commit_1_valid) begin
        if(_zz_134) begin
          rob_0_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_135) begin
          rob_1_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_136) begin
          rob_2_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_137) begin
          rob_3_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_138) begin
          rob_4_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_139) begin
          rob_5_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_140) begin
          rob_6_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_141) begin
          rob_7_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_142) begin
          rob_8_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_143) begin
          rob_9_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_144) begin
          rob_10_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_145) begin
          rob_11_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_146) begin
          rob_12_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_147) begin
          rob_13_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_148) begin
          rob_14_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_149) begin
          rob_15_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_150) begin
          rob_16_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_151) begin
          rob_17_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_152) begin
          rob_18_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_153) begin
          rob_19_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_154) begin
          rob_20_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_155) begin
          rob_21_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_156) begin
          rob_22_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_157) begin
          rob_23_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_158) begin
          rob_24_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_159) begin
          rob_25_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_160) begin
          rob_26_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_161) begin
          rob_27_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_162) begin
          rob_28_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_163) begin
          rob_29_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_164) begin
          rob_30_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_165) begin
          rob_31_branchResult_targetPC <= io_commit_1_branchResult_targetPC;
        end
        if(_zz_134) begin
          rob_0_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_135) begin
          rob_1_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_136) begin
          rob_2_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_137) begin
          rob_3_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_138) begin
          rob_4_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_139) begin
          rob_5_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_140) begin
          rob_6_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_141) begin
          rob_7_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_142) begin
          rob_8_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_143) begin
          rob_9_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_144) begin
          rob_10_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_145) begin
          rob_11_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_146) begin
          rob_12_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_147) begin
          rob_13_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_148) begin
          rob_14_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_149) begin
          rob_15_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_150) begin
          rob_16_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_151) begin
          rob_17_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_152) begin
          rob_18_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_153) begin
          rob_19_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_154) begin
          rob_20_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_155) begin
          rob_21_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_156) begin
          rob_22_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_157) begin
          rob_23_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_158) begin
          rob_24_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_159) begin
          rob_25_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_160) begin
          rob_26_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_161) begin
          rob_27_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_162) begin
          rob_28_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_163) begin
          rob_29_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_164) begin
          rob_30_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_165) begin
          rob_31_branchResult_branchResult <= io_commit_1_branchResult_branchResult;
        end
        if(_zz_134) begin
          rob_0_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_135) begin
          rob_1_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_136) begin
          rob_2_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_137) begin
          rob_3_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_138) begin
          rob_4_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_139) begin
          rob_5_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_140) begin
          rob_6_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_141) begin
          rob_7_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_142) begin
          rob_8_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_143) begin
          rob_9_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_144) begin
          rob_10_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_145) begin
          rob_11_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_146) begin
          rob_12_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_147) begin
          rob_13_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_148) begin
          rob_14_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_149) begin
          rob_15_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_150) begin
          rob_16_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_151) begin
          rob_17_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_152) begin
          rob_18_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_153) begin
          rob_19_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_154) begin
          rob_20_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_155) begin
          rob_21_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_156) begin
          rob_22_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_157) begin
          rob_23_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_158) begin
          rob_24_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_159) begin
          rob_25_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_160) begin
          rob_26_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_161) begin
          rob_27_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_162) begin
          rob_28_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_163) begin
          rob_29_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_164) begin
          rob_30_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_165) begin
          rob_31_branchResult_predictFail <= io_commit_1_branchResult_predictFail;
        end
        if(_zz_167) begin
          rob_0_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_168) begin
          rob_1_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_169) begin
          rob_2_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_170) begin
          rob_3_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_171) begin
          rob_4_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_172) begin
          rob_5_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_173) begin
          rob_6_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_174) begin
          rob_7_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_175) begin
          rob_8_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_176) begin
          rob_9_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_177) begin
          rob_10_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_178) begin
          rob_11_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_179) begin
          rob_12_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_180) begin
          rob_13_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_181) begin
          rob_14_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_182) begin
          rob_15_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_183) begin
          rob_16_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_184) begin
          rob_17_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_185) begin
          rob_18_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_186) begin
          rob_19_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_187) begin
          rob_20_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_188) begin
          rob_21_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_189) begin
          rob_22_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_190) begin
          rob_23_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_191) begin
          rob_24_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_192) begin
          rob_25_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_193) begin
          rob_26_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_194) begin
          rob_27_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_195) begin
          rob_28_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_196) begin
          rob_29_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_197) begin
          rob_30_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_198) begin
          rob_31_exceptionInfo_exception <= io_commit_1_exceptionInfo_exception;
        end
        if(_zz_167) begin
          rob_0_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_168) begin
          rob_1_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_169) begin
          rob_2_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_170) begin
          rob_3_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_171) begin
          rob_4_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_172) begin
          rob_5_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_173) begin
          rob_6_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_174) begin
          rob_7_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_175) begin
          rob_8_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_176) begin
          rob_9_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_177) begin
          rob_10_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_178) begin
          rob_11_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_179) begin
          rob_12_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_180) begin
          rob_13_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_181) begin
          rob_14_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_182) begin
          rob_15_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_183) begin
          rob_16_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_184) begin
          rob_17_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_185) begin
          rob_18_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_186) begin
          rob_19_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_187) begin
          rob_20_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_188) begin
          rob_21_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_189) begin
          rob_22_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_190) begin
          rob_23_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_191) begin
          rob_24_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_192) begin
          rob_25_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_193) begin
          rob_26_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_194) begin
          rob_27_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_195) begin
          rob_28_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_196) begin
          rob_29_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_197) begin
          rob_30_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_198) begin
          rob_31_exceptionInfo_eCode <= io_commit_1_exceptionInfo_eCode;
        end
        if(_zz_167) begin
          rob_0_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_168) begin
          rob_1_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_169) begin
          rob_2_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_170) begin
          rob_3_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_171) begin
          rob_4_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_172) begin
          rob_5_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_173) begin
          rob_6_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_174) begin
          rob_7_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_175) begin
          rob_8_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_176) begin
          rob_9_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_177) begin
          rob_10_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_178) begin
          rob_11_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_179) begin
          rob_12_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_180) begin
          rob_13_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_181) begin
          rob_14_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_182) begin
          rob_15_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_183) begin
          rob_16_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_184) begin
          rob_17_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_185) begin
          rob_18_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_186) begin
          rob_19_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_187) begin
          rob_20_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_188) begin
          rob_21_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_189) begin
          rob_22_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_190) begin
          rob_23_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_191) begin
          rob_24_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_192) begin
          rob_25_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_193) begin
          rob_26_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_194) begin
          rob_27_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_195) begin
          rob_28_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_196) begin
          rob_29_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_197) begin
          rob_30_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
        if(_zz_198) begin
          rob_31_exceptionInfo_eSubCode <= io_commit_1_exceptionInfo_eSubCode;
        end
      end
      if(io_commit_2_valid) begin
        if(_zz_200) begin
          rob_0_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_201) begin
          rob_1_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_202) begin
          rob_2_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_203) begin
          rob_3_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_204) begin
          rob_4_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_205) begin
          rob_5_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_206) begin
          rob_6_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_207) begin
          rob_7_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_208) begin
          rob_8_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_209) begin
          rob_9_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_210) begin
          rob_10_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_211) begin
          rob_11_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_212) begin
          rob_12_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_213) begin
          rob_13_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_214) begin
          rob_14_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_215) begin
          rob_15_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_216) begin
          rob_16_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_217) begin
          rob_17_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_218) begin
          rob_18_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_219) begin
          rob_19_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_220) begin
          rob_20_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_221) begin
          rob_21_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_222) begin
          rob_22_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_223) begin
          rob_23_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_224) begin
          rob_24_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_225) begin
          rob_25_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_226) begin
          rob_26_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_227) begin
          rob_27_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_228) begin
          rob_28_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_229) begin
          rob_29_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_230) begin
          rob_30_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_231) begin
          rob_31_branchResult_targetPC <= io_commit_2_branchResult_targetPC;
        end
        if(_zz_200) begin
          rob_0_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_201) begin
          rob_1_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_202) begin
          rob_2_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_203) begin
          rob_3_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_204) begin
          rob_4_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_205) begin
          rob_5_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_206) begin
          rob_6_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_207) begin
          rob_7_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_208) begin
          rob_8_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_209) begin
          rob_9_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_210) begin
          rob_10_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_211) begin
          rob_11_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_212) begin
          rob_12_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_213) begin
          rob_13_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_214) begin
          rob_14_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_215) begin
          rob_15_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_216) begin
          rob_16_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_217) begin
          rob_17_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_218) begin
          rob_18_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_219) begin
          rob_19_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_220) begin
          rob_20_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_221) begin
          rob_21_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_222) begin
          rob_22_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_223) begin
          rob_23_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_224) begin
          rob_24_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_225) begin
          rob_25_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_226) begin
          rob_26_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_227) begin
          rob_27_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_228) begin
          rob_28_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_229) begin
          rob_29_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_230) begin
          rob_30_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_231) begin
          rob_31_branchResult_branchResult <= io_commit_2_branchResult_branchResult;
        end
        if(_zz_200) begin
          rob_0_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_201) begin
          rob_1_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_202) begin
          rob_2_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_203) begin
          rob_3_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_204) begin
          rob_4_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_205) begin
          rob_5_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_206) begin
          rob_6_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_207) begin
          rob_7_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_208) begin
          rob_8_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_209) begin
          rob_9_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_210) begin
          rob_10_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_211) begin
          rob_11_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_212) begin
          rob_12_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_213) begin
          rob_13_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_214) begin
          rob_14_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_215) begin
          rob_15_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_216) begin
          rob_16_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_217) begin
          rob_17_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_218) begin
          rob_18_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_219) begin
          rob_19_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_220) begin
          rob_20_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_221) begin
          rob_21_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_222) begin
          rob_22_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_223) begin
          rob_23_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_224) begin
          rob_24_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_225) begin
          rob_25_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_226) begin
          rob_26_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_227) begin
          rob_27_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_228) begin
          rob_28_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_229) begin
          rob_29_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_230) begin
          rob_30_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_231) begin
          rob_31_branchResult_predictFail <= io_commit_2_branchResult_predictFail;
        end
        if(_zz_233) begin
          rob_0_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_234) begin
          rob_1_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_235) begin
          rob_2_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_236) begin
          rob_3_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_237) begin
          rob_4_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_238) begin
          rob_5_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_239) begin
          rob_6_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_240) begin
          rob_7_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_241) begin
          rob_8_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_242) begin
          rob_9_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_243) begin
          rob_10_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_244) begin
          rob_11_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_245) begin
          rob_12_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_246) begin
          rob_13_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_247) begin
          rob_14_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_248) begin
          rob_15_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_249) begin
          rob_16_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_250) begin
          rob_17_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_251) begin
          rob_18_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_252) begin
          rob_19_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_253) begin
          rob_20_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_254) begin
          rob_21_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_255) begin
          rob_22_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_256) begin
          rob_23_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_257) begin
          rob_24_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_258) begin
          rob_25_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_259) begin
          rob_26_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_260) begin
          rob_27_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_261) begin
          rob_28_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_262) begin
          rob_29_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_263) begin
          rob_30_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_264) begin
          rob_31_exceptionInfo_exception <= io_commit_2_exceptionInfo_exception;
        end
        if(_zz_233) begin
          rob_0_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_234) begin
          rob_1_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_235) begin
          rob_2_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_236) begin
          rob_3_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_237) begin
          rob_4_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_238) begin
          rob_5_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_239) begin
          rob_6_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_240) begin
          rob_7_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_241) begin
          rob_8_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_242) begin
          rob_9_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_243) begin
          rob_10_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_244) begin
          rob_11_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_245) begin
          rob_12_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_246) begin
          rob_13_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_247) begin
          rob_14_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_248) begin
          rob_15_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_249) begin
          rob_16_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_250) begin
          rob_17_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_251) begin
          rob_18_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_252) begin
          rob_19_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_253) begin
          rob_20_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_254) begin
          rob_21_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_255) begin
          rob_22_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_256) begin
          rob_23_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_257) begin
          rob_24_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_258) begin
          rob_25_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_259) begin
          rob_26_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_260) begin
          rob_27_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_261) begin
          rob_28_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_262) begin
          rob_29_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_263) begin
          rob_30_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_264) begin
          rob_31_exceptionInfo_eCode <= io_commit_2_exceptionInfo_eCode;
        end
        if(_zz_233) begin
          rob_0_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_234) begin
          rob_1_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_235) begin
          rob_2_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_236) begin
          rob_3_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_237) begin
          rob_4_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_238) begin
          rob_5_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_239) begin
          rob_6_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_240) begin
          rob_7_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_241) begin
          rob_8_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_242) begin
          rob_9_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_243) begin
          rob_10_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_244) begin
          rob_11_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_245) begin
          rob_12_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_246) begin
          rob_13_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_247) begin
          rob_14_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_248) begin
          rob_15_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_249) begin
          rob_16_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_250) begin
          rob_17_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_251) begin
          rob_18_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_252) begin
          rob_19_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_253) begin
          rob_20_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_254) begin
          rob_21_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_255) begin
          rob_22_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_256) begin
          rob_23_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_257) begin
          rob_24_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_258) begin
          rob_25_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_259) begin
          rob_26_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_260) begin
          rob_27_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_261) begin
          rob_28_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_262) begin
          rob_29_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_263) begin
          rob_30_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
        if(_zz_264) begin
          rob_31_exceptionInfo_eSubCode <= io_commit_2_exceptionInfo_eSubCode;
        end
      end
      if(io_commit_3_valid) begin
        if(_zz_266) begin
          rob_0_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_267) begin
          rob_1_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_268) begin
          rob_2_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_269) begin
          rob_3_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_270) begin
          rob_4_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_271) begin
          rob_5_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_272) begin
          rob_6_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_273) begin
          rob_7_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_274) begin
          rob_8_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_275) begin
          rob_9_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_276) begin
          rob_10_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_277) begin
          rob_11_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_278) begin
          rob_12_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_279) begin
          rob_13_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_280) begin
          rob_14_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_281) begin
          rob_15_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_282) begin
          rob_16_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_283) begin
          rob_17_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_284) begin
          rob_18_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_285) begin
          rob_19_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_286) begin
          rob_20_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_287) begin
          rob_21_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_288) begin
          rob_22_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_289) begin
          rob_23_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_290) begin
          rob_24_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_291) begin
          rob_25_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_292) begin
          rob_26_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_293) begin
          rob_27_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_294) begin
          rob_28_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_295) begin
          rob_29_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_296) begin
          rob_30_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_297) begin
          rob_31_branchResult_targetPC <= io_commit_3_branchResult_targetPC;
        end
        if(_zz_266) begin
          rob_0_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_267) begin
          rob_1_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_268) begin
          rob_2_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_269) begin
          rob_3_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_270) begin
          rob_4_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_271) begin
          rob_5_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_272) begin
          rob_6_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_273) begin
          rob_7_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_274) begin
          rob_8_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_275) begin
          rob_9_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_276) begin
          rob_10_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_277) begin
          rob_11_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_278) begin
          rob_12_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_279) begin
          rob_13_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_280) begin
          rob_14_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_281) begin
          rob_15_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_282) begin
          rob_16_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_283) begin
          rob_17_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_284) begin
          rob_18_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_285) begin
          rob_19_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_286) begin
          rob_20_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_287) begin
          rob_21_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_288) begin
          rob_22_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_289) begin
          rob_23_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_290) begin
          rob_24_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_291) begin
          rob_25_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_292) begin
          rob_26_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_293) begin
          rob_27_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_294) begin
          rob_28_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_295) begin
          rob_29_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_296) begin
          rob_30_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_297) begin
          rob_31_branchResult_branchResult <= io_commit_3_branchResult_branchResult;
        end
        if(_zz_266) begin
          rob_0_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_267) begin
          rob_1_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_268) begin
          rob_2_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_269) begin
          rob_3_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_270) begin
          rob_4_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_271) begin
          rob_5_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_272) begin
          rob_6_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_273) begin
          rob_7_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_274) begin
          rob_8_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_275) begin
          rob_9_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_276) begin
          rob_10_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_277) begin
          rob_11_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_278) begin
          rob_12_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_279) begin
          rob_13_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_280) begin
          rob_14_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_281) begin
          rob_15_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_282) begin
          rob_16_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_283) begin
          rob_17_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_284) begin
          rob_18_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_285) begin
          rob_19_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_286) begin
          rob_20_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_287) begin
          rob_21_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_288) begin
          rob_22_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_289) begin
          rob_23_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_290) begin
          rob_24_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_291) begin
          rob_25_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_292) begin
          rob_26_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_293) begin
          rob_27_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_294) begin
          rob_28_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_295) begin
          rob_29_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_296) begin
          rob_30_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_297) begin
          rob_31_branchResult_predictFail <= io_commit_3_branchResult_predictFail;
        end
        if(_zz_299) begin
          rob_0_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_300) begin
          rob_1_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_301) begin
          rob_2_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_302) begin
          rob_3_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_303) begin
          rob_4_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_304) begin
          rob_5_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_305) begin
          rob_6_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_306) begin
          rob_7_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_307) begin
          rob_8_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_308) begin
          rob_9_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_309) begin
          rob_10_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_310) begin
          rob_11_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_311) begin
          rob_12_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_312) begin
          rob_13_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_313) begin
          rob_14_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_314) begin
          rob_15_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_315) begin
          rob_16_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_316) begin
          rob_17_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_317) begin
          rob_18_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_318) begin
          rob_19_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_319) begin
          rob_20_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_320) begin
          rob_21_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_321) begin
          rob_22_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_322) begin
          rob_23_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_323) begin
          rob_24_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_324) begin
          rob_25_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_325) begin
          rob_26_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_326) begin
          rob_27_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_327) begin
          rob_28_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_328) begin
          rob_29_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_329) begin
          rob_30_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_330) begin
          rob_31_exceptionInfo_exception <= io_commit_3_exceptionInfo_exception;
        end
        if(_zz_299) begin
          rob_0_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_300) begin
          rob_1_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_301) begin
          rob_2_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_302) begin
          rob_3_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_303) begin
          rob_4_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_304) begin
          rob_5_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_305) begin
          rob_6_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_306) begin
          rob_7_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_307) begin
          rob_8_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_308) begin
          rob_9_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_309) begin
          rob_10_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_310) begin
          rob_11_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_311) begin
          rob_12_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_312) begin
          rob_13_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_313) begin
          rob_14_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_314) begin
          rob_15_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_315) begin
          rob_16_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_316) begin
          rob_17_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_317) begin
          rob_18_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_318) begin
          rob_19_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_319) begin
          rob_20_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_320) begin
          rob_21_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_321) begin
          rob_22_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_322) begin
          rob_23_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_323) begin
          rob_24_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_324) begin
          rob_25_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_325) begin
          rob_26_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_326) begin
          rob_27_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_327) begin
          rob_28_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_328) begin
          rob_29_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_329) begin
          rob_30_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_330) begin
          rob_31_exceptionInfo_eCode <= io_commit_3_exceptionInfo_eCode;
        end
        if(_zz_299) begin
          rob_0_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_300) begin
          rob_1_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_301) begin
          rob_2_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_302) begin
          rob_3_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_303) begin
          rob_4_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_304) begin
          rob_5_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_305) begin
          rob_6_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_306) begin
          rob_7_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_307) begin
          rob_8_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_308) begin
          rob_9_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_309) begin
          rob_10_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_310) begin
          rob_11_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_311) begin
          rob_12_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_312) begin
          rob_13_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_313) begin
          rob_14_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_314) begin
          rob_15_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_315) begin
          rob_16_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_316) begin
          rob_17_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_317) begin
          rob_18_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_318) begin
          rob_19_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_319) begin
          rob_20_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_320) begin
          rob_21_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_321) begin
          rob_22_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_322) begin
          rob_23_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_323) begin
          rob_24_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_324) begin
          rob_25_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_325) begin
          rob_26_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_326) begin
          rob_27_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_327) begin
          rob_28_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_328) begin
          rob_29_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_329) begin
          rob_30_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
        if(_zz_330) begin
          rob_31_exceptionInfo_eSubCode <= io_commit_3_exceptionInfo_eSubCode;
        end
      end
      if(io_commit_4_valid) begin
        if(_zz_332) begin
          rob_0_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_333) begin
          rob_1_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_334) begin
          rob_2_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_335) begin
          rob_3_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_336) begin
          rob_4_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_337) begin
          rob_5_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_338) begin
          rob_6_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_339) begin
          rob_7_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_340) begin
          rob_8_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_341) begin
          rob_9_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_342) begin
          rob_10_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_343) begin
          rob_11_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_344) begin
          rob_12_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_345) begin
          rob_13_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_346) begin
          rob_14_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_347) begin
          rob_15_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_348) begin
          rob_16_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_349) begin
          rob_17_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_350) begin
          rob_18_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_351) begin
          rob_19_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_352) begin
          rob_20_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_353) begin
          rob_21_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_354) begin
          rob_22_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_355) begin
          rob_23_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_356) begin
          rob_24_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_357) begin
          rob_25_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_358) begin
          rob_26_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_359) begin
          rob_27_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_360) begin
          rob_28_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_361) begin
          rob_29_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_362) begin
          rob_30_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_363) begin
          rob_31_branchResult_targetPC <= io_commit_4_branchResult_targetPC;
        end
        if(_zz_332) begin
          rob_0_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_333) begin
          rob_1_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_334) begin
          rob_2_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_335) begin
          rob_3_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_336) begin
          rob_4_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_337) begin
          rob_5_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_338) begin
          rob_6_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_339) begin
          rob_7_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_340) begin
          rob_8_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_341) begin
          rob_9_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_342) begin
          rob_10_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_343) begin
          rob_11_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_344) begin
          rob_12_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_345) begin
          rob_13_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_346) begin
          rob_14_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_347) begin
          rob_15_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_348) begin
          rob_16_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_349) begin
          rob_17_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_350) begin
          rob_18_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_351) begin
          rob_19_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_352) begin
          rob_20_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_353) begin
          rob_21_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_354) begin
          rob_22_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_355) begin
          rob_23_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_356) begin
          rob_24_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_357) begin
          rob_25_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_358) begin
          rob_26_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_359) begin
          rob_27_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_360) begin
          rob_28_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_361) begin
          rob_29_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_362) begin
          rob_30_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_363) begin
          rob_31_branchResult_branchResult <= io_commit_4_branchResult_branchResult;
        end
        if(_zz_332) begin
          rob_0_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_333) begin
          rob_1_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_334) begin
          rob_2_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_335) begin
          rob_3_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_336) begin
          rob_4_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_337) begin
          rob_5_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_338) begin
          rob_6_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_339) begin
          rob_7_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_340) begin
          rob_8_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_341) begin
          rob_9_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_342) begin
          rob_10_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_343) begin
          rob_11_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_344) begin
          rob_12_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_345) begin
          rob_13_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_346) begin
          rob_14_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_347) begin
          rob_15_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_348) begin
          rob_16_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_349) begin
          rob_17_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_350) begin
          rob_18_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_351) begin
          rob_19_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_352) begin
          rob_20_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_353) begin
          rob_21_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_354) begin
          rob_22_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_355) begin
          rob_23_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_356) begin
          rob_24_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_357) begin
          rob_25_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_358) begin
          rob_26_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_359) begin
          rob_27_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_360) begin
          rob_28_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_361) begin
          rob_29_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_362) begin
          rob_30_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_363) begin
          rob_31_branchResult_predictFail <= io_commit_4_branchResult_predictFail;
        end
        if(_zz_365) begin
          rob_0_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_366) begin
          rob_1_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_367) begin
          rob_2_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_368) begin
          rob_3_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_369) begin
          rob_4_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_370) begin
          rob_5_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_371) begin
          rob_6_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_372) begin
          rob_7_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_373) begin
          rob_8_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_374) begin
          rob_9_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_375) begin
          rob_10_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_376) begin
          rob_11_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_377) begin
          rob_12_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_378) begin
          rob_13_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_379) begin
          rob_14_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_380) begin
          rob_15_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_381) begin
          rob_16_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_382) begin
          rob_17_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_383) begin
          rob_18_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_384) begin
          rob_19_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_385) begin
          rob_20_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_386) begin
          rob_21_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_387) begin
          rob_22_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_388) begin
          rob_23_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_389) begin
          rob_24_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_390) begin
          rob_25_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_391) begin
          rob_26_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_392) begin
          rob_27_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_393) begin
          rob_28_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_394) begin
          rob_29_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_395) begin
          rob_30_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_396) begin
          rob_31_exceptionInfo_exception <= io_commit_4_exceptionInfo_exception;
        end
        if(_zz_365) begin
          rob_0_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_366) begin
          rob_1_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_367) begin
          rob_2_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_368) begin
          rob_3_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_369) begin
          rob_4_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_370) begin
          rob_5_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_371) begin
          rob_6_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_372) begin
          rob_7_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_373) begin
          rob_8_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_374) begin
          rob_9_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_375) begin
          rob_10_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_376) begin
          rob_11_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_377) begin
          rob_12_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_378) begin
          rob_13_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_379) begin
          rob_14_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_380) begin
          rob_15_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_381) begin
          rob_16_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_382) begin
          rob_17_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_383) begin
          rob_18_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_384) begin
          rob_19_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_385) begin
          rob_20_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_386) begin
          rob_21_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_387) begin
          rob_22_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_388) begin
          rob_23_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_389) begin
          rob_24_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_390) begin
          rob_25_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_391) begin
          rob_26_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_392) begin
          rob_27_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_393) begin
          rob_28_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_394) begin
          rob_29_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_395) begin
          rob_30_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_396) begin
          rob_31_exceptionInfo_eCode <= io_commit_4_exceptionInfo_eCode;
        end
        if(_zz_365) begin
          rob_0_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_366) begin
          rob_1_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_367) begin
          rob_2_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_368) begin
          rob_3_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_369) begin
          rob_4_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_370) begin
          rob_5_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_371) begin
          rob_6_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_372) begin
          rob_7_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_373) begin
          rob_8_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_374) begin
          rob_9_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_375) begin
          rob_10_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_376) begin
          rob_11_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_377) begin
          rob_12_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_378) begin
          rob_13_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_379) begin
          rob_14_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_380) begin
          rob_15_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_381) begin
          rob_16_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_382) begin
          rob_17_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_383) begin
          rob_18_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_384) begin
          rob_19_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_385) begin
          rob_20_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_386) begin
          rob_21_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_387) begin
          rob_22_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_388) begin
          rob_23_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_389) begin
          rob_24_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_390) begin
          rob_25_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_391) begin
          rob_26_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_392) begin
          rob_27_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_393) begin
          rob_28_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_394) begin
          rob_29_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_395) begin
          rob_30_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
        if(_zz_396) begin
          rob_31_exceptionInfo_eSubCode <= io_commit_4_exceptionInfo_eSubCode;
        end
      end
      head_0 <= (io_flush ? 5'h00 : _zz_head_0);
      head_1 <= (io_flush ? 5'h01 : _zz_head_1);
      delayedFlush <= io_flush;
      stageReg_availROBMask <= (io_flush ? 2'b00 : stage_availROBMask);
      stageReg_retireARAT_0_ard <= (io_flush ? 5'h00 : stage_retireARAT_0_ard);
      stageReg_retireARAT_0_prd <= (io_flush ? 6'h00 : stage_retireARAT_0_prd);
      stageReg_retireARAT_0_wen <= (io_flush ? 1'b0 : stage_retireARAT_0_wen);
      stageReg_retireARAT_1_ard <= (io_flush ? 5'h00 : stage_retireARAT_1_ard);
      stageReg_retireARAT_1_prd <= (io_flush ? 6'h00 : stage_retireARAT_1_prd);
      stageReg_retireARAT_1_wen <= (io_flush ? 1'b0 : stage_retireARAT_1_wen);
      stageReg_freePRFIdx_0 <= (io_flush ? 6'h00 : stage_freePRFIdx_0);
      stageReg_freePRFIdx_1 <= (io_flush ? 6'h00 : stage_freePRFIdx_1);
      stageReg_freePRFNum <= (io_flush ? 2'b00 : stage_freePRFNum);
      stageReg_retireROBIdx_0 <= (io_flush ? 5'h00 : stage_retireROBIdx_0);
      stageReg_retireROBIdx_1 <= (io_flush ? 5'h00 : stage_retireROBIdx_1);
      stageReg_retireEn_0 <= (io_flush ? 1'b0 : stage_retireEn_0);
      stageReg_retireEn_1 <= (io_flush ? 1'b0 : stage_retireEn_1);
      stageReg_wakeupMem <= (io_flush ? 1'b0 : stage_wakeupMem);
      stageReg_retireLLBitUpdate <= (io_flush ? 1'b0 : stage_retireLLBitUpdate);
      stageReg_retireWriteCSR <= (io_flush ? 1'b0 : stage_retireWriteCSR);
      stageReg_retireERTN <= (io_flush ? 1'b0 : stage_retireERTN);
      stageReg_retireNormalException <= (io_flush ? 1'b0 : stage_retireNormalException);
      stageReg_retireTLBRException <= (io_flush ? 1'b0 : stage_retireTLBRException);
      stageReg_retireEPC <= (io_flush ? 32'h00000000 : stage_retireEPC);
      stageReg_retireEROBIdx <= (io_flush ? 5'h00 : stage_retireEROBIdx);
      stageReg_retireECode <= (io_flush ? 6'h00 : stage_retireECode);
      stageReg_retireESubCode <= (io_flush ? 1'b0 : stage_retireESubCode);
      stageReg_updateBPU_0_pc <= (io_flush ? 32'h00000000 : stage_updateBPU_0_pc);
      stageReg_updateBPU_0_isJumpInst <= (io_flush ? 1'b0 : stage_updateBPU_0_isJumpInst);
      stageReg_updateBPU_0_taken <= (io_flush ? 1'b0 : stage_updateBPU_0_taken);
      stageReg_updateBPU_0_predictFail <= (io_flush ? 1'b0 : stage_updateBPU_0_predictFail);
      stageReg_updateBPU_0_target <= (io_flush ? 32'h00000000 : stage_updateBPU_0_target);
      stageReg_updateBPU_1_pc <= (io_flush ? 32'h00000000 : stage_updateBPU_1_pc);
      stageReg_updateBPU_1_isJumpInst <= (io_flush ? 1'b0 : stage_updateBPU_1_isJumpInst);
      stageReg_updateBPU_1_taken <= (io_flush ? 1'b0 : stage_updateBPU_1_taken);
      stageReg_updateBPU_1_predictFail <= (io_flush ? 1'b0 : stage_updateBPU_1_predictFail);
      stageReg_updateBPU_1_target <= (io_flush ? 32'h00000000 : stage_updateBPU_1_target);
      stageReg_flush <= (io_flush ? 1'b0 : stage_flush);
      stageReg_redirectPC <= (io_flush ? 32'h00000000 : stage_redirectPC);
    end
  end


endmodule

module PRF (
  input  wire [5:0]    io_read_0_0_idx,
  output reg  [31:0]   io_read_0_0_data,
  input  wire [5:0]    io_read_0_1_idx,
  output reg  [31:0]   io_read_0_1_data,
  input  wire [5:0]    io_read_1_0_idx,
  output reg  [31:0]   io_read_1_0_data,
  input  wire [5:0]    io_read_1_1_idx,
  output reg  [31:0]   io_read_1_1_data,
  input  wire [5:0]    io_read_2_0_idx,
  output reg  [31:0]   io_read_2_0_data,
  input  wire [5:0]    io_read_2_1_idx,
  output reg  [31:0]   io_read_2_1_data,
  input  wire [5:0]    io_read_3_0_idx,
  output reg  [31:0]   io_read_3_0_data,
  input  wire [5:0]    io_read_3_1_idx,
  output reg  [31:0]   io_read_3_1_data,
  input  wire [5:0]    io_read_4_0_idx,
  output reg  [31:0]   io_read_4_0_data,
  input  wire [5:0]    io_read_4_1_idx,
  output reg  [31:0]   io_read_4_1_data,
  input  wire [5:0]    io_write_0_idx,
  input  wire [31:0]   io_write_0_data,
  input  wire [5:0]    io_write_1_idx,
  input  wire [31:0]   io_write_1_data,
  input  wire [5:0]    io_write_2_idx,
  input  wire [31:0]   io_write_2_data,
  input  wire [5:0]    io_write_3_idx,
  input  wire [31:0]   io_write_3_data,
  input  wire [5:0]    io_write_4_idx,
  input  wire [31:0]   io_write_4_data,
  output reg  [31:0]   io_debugRegs_0,
  output reg  [31:0]   io_debugRegs_1,
  output reg  [31:0]   io_debugRegs_2,
  output reg  [31:0]   io_debugRegs_3,
  output reg  [31:0]   io_debugRegs_4,
  output reg  [31:0]   io_debugRegs_5,
  output reg  [31:0]   io_debugRegs_6,
  output reg  [31:0]   io_debugRegs_7,
  output reg  [31:0]   io_debugRegs_8,
  output reg  [31:0]   io_debugRegs_9,
  output reg  [31:0]   io_debugRegs_10,
  output reg  [31:0]   io_debugRegs_11,
  output reg  [31:0]   io_debugRegs_12,
  output reg  [31:0]   io_debugRegs_13,
  output reg  [31:0]   io_debugRegs_14,
  output reg  [31:0]   io_debugRegs_15,
  output reg  [31:0]   io_debugRegs_16,
  output reg  [31:0]   io_debugRegs_17,
  output reg  [31:0]   io_debugRegs_18,
  output reg  [31:0]   io_debugRegs_19,
  output reg  [31:0]   io_debugRegs_20,
  output reg  [31:0]   io_debugRegs_21,
  output reg  [31:0]   io_debugRegs_22,
  output reg  [31:0]   io_debugRegs_23,
  output reg  [31:0]   io_debugRegs_24,
  output reg  [31:0]   io_debugRegs_25,
  output reg  [31:0]   io_debugRegs_26,
  output reg  [31:0]   io_debugRegs_27,
  output reg  [31:0]   io_debugRegs_28,
  output reg  [31:0]   io_debugRegs_29,
  output reg  [31:0]   io_debugRegs_30,
  output reg  [31:0]   io_debugRegs_31,
  output reg  [31:0]   io_debugRegs_32,
  output reg  [31:0]   io_debugRegs_33,
  output reg  [31:0]   io_debugRegs_34,
  output reg  [31:0]   io_debugRegs_35,
  output reg  [31:0]   io_debugRegs_36,
  output reg  [31:0]   io_debugRegs_37,
  output reg  [31:0]   io_debugRegs_38,
  output reg  [31:0]   io_debugRegs_39,
  output reg  [31:0]   io_debugRegs_40,
  output reg  [31:0]   io_debugRegs_41,
  output reg  [31:0]   io_debugRegs_42,
  output reg  [31:0]   io_debugRegs_43,
  output reg  [31:0]   io_debugRegs_44,
  output reg  [31:0]   io_debugRegs_45,
  output reg  [31:0]   io_debugRegs_46,
  output reg  [31:0]   io_debugRegs_47,
  output reg  [31:0]   io_debugRegs_48,
  output reg  [31:0]   io_debugRegs_49,
  output reg  [31:0]   io_debugRegs_50,
  output reg  [31:0]   io_debugRegs_51,
  output reg  [31:0]   io_debugRegs_52,
  output reg  [31:0]   io_debugRegs_53,
  output reg  [31:0]   io_debugRegs_54,
  output reg  [31:0]   io_debugRegs_55,
  output reg  [31:0]   io_debugRegs_56,
  output reg  [31:0]   io_debugRegs_57,
  output reg  [31:0]   io_debugRegs_58,
  output reg  [31:0]   io_debugRegs_59,
  output reg  [31:0]   io_debugRegs_60,
  output reg  [31:0]   io_debugRegs_61,
  output reg  [31:0]   io_debugRegs_62,
  output reg  [31:0]   io_debugRegs_63,
  input  wire          aclk,
  input  wire          aresetn
);

  wire       [5:0]    _zz_when_PRF_l19;
  wire       [0:0]    _zz_when_PRF_l19_1;
  reg        [31:0]   _zz_io_read_0_0_data;
  wire       [5:0]    _zz_io_read_0_0_data_1;
  wire       [0:0]    _zz_io_read_0_0_data_2;
  wire       [5:0]    _zz_when_PRF_l19_1_1;
  wire       [0:0]    _zz_when_PRF_l19_1_2;
  reg        [31:0]   _zz_io_read_0_1_data;
  wire       [5:0]    _zz_io_read_0_1_data_1;
  wire       [0:0]    _zz_io_read_0_1_data_2;
  wire       [5:0]    _zz_when_PRF_l19_2;
  wire       [0:0]    _zz_when_PRF_l19_2_1;
  reg        [31:0]   _zz_io_read_1_0_data;
  wire       [5:0]    _zz_io_read_1_0_data_1;
  wire       [0:0]    _zz_io_read_1_0_data_2;
  wire       [5:0]    _zz_when_PRF_l19_3;
  wire       [0:0]    _zz_when_PRF_l19_3_1;
  reg        [31:0]   _zz_io_read_1_1_data;
  wire       [5:0]    _zz_io_read_1_1_data_1;
  wire       [0:0]    _zz_io_read_1_1_data_2;
  wire       [5:0]    _zz_when_PRF_l19_4;
  wire       [0:0]    _zz_when_PRF_l19_4_1;
  reg        [31:0]   _zz_io_read_2_0_data;
  wire       [5:0]    _zz_io_read_2_0_data_1;
  wire       [0:0]    _zz_io_read_2_0_data_2;
  wire       [5:0]    _zz_when_PRF_l19_5;
  wire       [0:0]    _zz_when_PRF_l19_5_1;
  reg        [31:0]   _zz_io_read_2_1_data;
  wire       [5:0]    _zz_io_read_2_1_data_1;
  wire       [0:0]    _zz_io_read_2_1_data_2;
  wire       [5:0]    _zz_when_PRF_l19_6;
  wire       [0:0]    _zz_when_PRF_l19_6_1;
  reg        [31:0]   _zz_io_read_3_0_data;
  wire       [5:0]    _zz_io_read_3_0_data_1;
  wire       [0:0]    _zz_io_read_3_0_data_2;
  wire       [5:0]    _zz_when_PRF_l19_7;
  wire       [0:0]    _zz_when_PRF_l19_7_1;
  reg        [31:0]   _zz_io_read_3_1_data;
  wire       [5:0]    _zz_io_read_3_1_data_1;
  wire       [0:0]    _zz_io_read_3_1_data_2;
  wire       [5:0]    _zz_when_PRF_l19_8;
  wire       [0:0]    _zz_when_PRF_l19_8_1;
  reg        [31:0]   _zz_io_read_4_0_data;
  wire       [5:0]    _zz_io_read_4_0_data_1;
  wire       [0:0]    _zz_io_read_4_0_data_2;
  wire       [5:0]    _zz_when_PRF_l19_9;
  wire       [0:0]    _zz_when_PRF_l19_9_1;
  reg        [31:0]   _zz_io_read_4_1_data;
  wire       [5:0]    _zz_io_read_4_1_data_1;
  wire       [0:0]    _zz_io_read_4_1_data_2;
  wire       [5:0]    _zz_when_PRF_l27;
  wire       [0:0]    _zz_when_PRF_l27_1;
  wire       [5:0]    _zz_when_PRF_l27_1_1;
  wire       [0:0]    _zz_when_PRF_l27_1_2;
  wire       [5:0]    _zz_when_PRF_l27_2;
  wire       [0:0]    _zz_when_PRF_l27_2_1;
  wire       [5:0]    _zz_when_PRF_l27_3;
  wire       [0:0]    _zz_when_PRF_l27_3_1;
  wire       [5:0]    _zz_when_PRF_l27_4;
  wire       [0:0]    _zz_when_PRF_l27_4_1;
  reg        [31:0]   regFile_0;
  reg        [31:0]   regFile_1;
  reg        [31:0]   regFile_2;
  reg        [31:0]   regFile_3;
  reg        [31:0]   regFile_4;
  reg        [31:0]   regFile_5;
  reg        [31:0]   regFile_6;
  reg        [31:0]   regFile_7;
  reg        [31:0]   regFile_8;
  reg        [31:0]   regFile_9;
  reg        [31:0]   regFile_10;
  reg        [31:0]   regFile_11;
  reg        [31:0]   regFile_12;
  reg        [31:0]   regFile_13;
  reg        [31:0]   regFile_14;
  reg        [31:0]   regFile_15;
  reg        [31:0]   regFile_16;
  reg        [31:0]   regFile_17;
  reg        [31:0]   regFile_18;
  reg        [31:0]   regFile_19;
  reg        [31:0]   regFile_20;
  reg        [31:0]   regFile_21;
  reg        [31:0]   regFile_22;
  reg        [31:0]   regFile_23;
  reg        [31:0]   regFile_24;
  reg        [31:0]   regFile_25;
  reg        [31:0]   regFile_26;
  reg        [31:0]   regFile_27;
  reg        [31:0]   regFile_28;
  reg        [31:0]   regFile_29;
  reg        [31:0]   regFile_30;
  reg        [31:0]   regFile_31;
  reg        [31:0]   regFile_32;
  reg        [31:0]   regFile_33;
  reg        [31:0]   regFile_34;
  reg        [31:0]   regFile_35;
  reg        [31:0]   regFile_36;
  reg        [31:0]   regFile_37;
  reg        [31:0]   regFile_38;
  reg        [31:0]   regFile_39;
  reg        [31:0]   regFile_40;
  reg        [31:0]   regFile_41;
  reg        [31:0]   regFile_42;
  reg        [31:0]   regFile_43;
  reg        [31:0]   regFile_44;
  reg        [31:0]   regFile_45;
  reg        [31:0]   regFile_46;
  reg        [31:0]   regFile_47;
  reg        [31:0]   regFile_48;
  reg        [31:0]   regFile_49;
  reg        [31:0]   regFile_50;
  reg        [31:0]   regFile_51;
  reg        [31:0]   regFile_52;
  reg        [31:0]   regFile_53;
  reg        [31:0]   regFile_54;
  reg        [31:0]   regFile_55;
  reg        [31:0]   regFile_56;
  reg        [31:0]   regFile_57;
  reg        [31:0]   regFile_58;
  reg        [31:0]   regFile_59;
  reg        [31:0]   regFile_60;
  reg        [31:0]   regFile_61;
  reg        [31:0]   regFile_62;
  reg        [31:0]   regFile_63;
  wire                when_PRF_l19;
  wire                when_PRF_l19_1;
  wire                when_PRF_l19_2;
  wire                when_PRF_l19_3;
  wire                when_PRF_l19_4;
  wire                when_PRF_l19_5;
  wire                when_PRF_l19_6;
  wire                when_PRF_l19_7;
  wire                when_PRF_l19_8;
  wire                when_PRF_l19_9;
  wire                when_PRF_l27;
  wire       [63:0]   _zz_1;
  wire                when_PRF_l27_1;
  wire       [63:0]   _zz_2;
  wire                when_PRF_l27_2;
  wire       [63:0]   _zz_3;
  wire                when_PRF_l27_3;
  wire       [63:0]   _zz_4;
  wire                when_PRF_l27_4;
  wire       [63:0]   _zz_5;

  assign _zz_when_PRF_l19_1 = 1'b0;
  assign _zz_when_PRF_l19 = {5'd0, _zz_when_PRF_l19_1};
  assign _zz_io_read_0_0_data_2 = 1'b0;
  assign _zz_when_PRF_l19_1_2 = 1'b0;
  assign _zz_when_PRF_l19_1_1 = {5'd0, _zz_when_PRF_l19_1_2};
  assign _zz_io_read_0_1_data_2 = 1'b0;
  assign _zz_when_PRF_l19_2_1 = 1'b0;
  assign _zz_when_PRF_l19_2 = {5'd0, _zz_when_PRF_l19_2_1};
  assign _zz_io_read_1_0_data_2 = 1'b0;
  assign _zz_when_PRF_l19_3_1 = 1'b0;
  assign _zz_when_PRF_l19_3 = {5'd0, _zz_when_PRF_l19_3_1};
  assign _zz_io_read_1_1_data_2 = 1'b0;
  assign _zz_when_PRF_l19_4_1 = 1'b0;
  assign _zz_when_PRF_l19_4 = {5'd0, _zz_when_PRF_l19_4_1};
  assign _zz_io_read_2_0_data_2 = 1'b0;
  assign _zz_when_PRF_l19_5_1 = 1'b0;
  assign _zz_when_PRF_l19_5 = {5'd0, _zz_when_PRF_l19_5_1};
  assign _zz_io_read_2_1_data_2 = 1'b0;
  assign _zz_when_PRF_l19_6_1 = 1'b0;
  assign _zz_when_PRF_l19_6 = {5'd0, _zz_when_PRF_l19_6_1};
  assign _zz_io_read_3_0_data_2 = 1'b0;
  assign _zz_when_PRF_l19_7_1 = 1'b0;
  assign _zz_when_PRF_l19_7 = {5'd0, _zz_when_PRF_l19_7_1};
  assign _zz_io_read_3_1_data_2 = 1'b0;
  assign _zz_when_PRF_l19_8_1 = 1'b0;
  assign _zz_when_PRF_l19_8 = {5'd0, _zz_when_PRF_l19_8_1};
  assign _zz_io_read_4_0_data_2 = 1'b0;
  assign _zz_when_PRF_l19_9_1 = 1'b0;
  assign _zz_when_PRF_l19_9 = {5'd0, _zz_when_PRF_l19_9_1};
  assign _zz_io_read_4_1_data_2 = 1'b0;
  assign _zz_when_PRF_l27_1 = 1'b0;
  assign _zz_when_PRF_l27 = {5'd0, _zz_when_PRF_l27_1};
  assign _zz_when_PRF_l27_1_2 = 1'b0;
  assign _zz_when_PRF_l27_1_1 = {5'd0, _zz_when_PRF_l27_1_2};
  assign _zz_when_PRF_l27_2_1 = 1'b0;
  assign _zz_when_PRF_l27_2 = {5'd0, _zz_when_PRF_l27_2_1};
  assign _zz_when_PRF_l27_3_1 = 1'b0;
  assign _zz_when_PRF_l27_3 = {5'd0, _zz_when_PRF_l27_3_1};
  assign _zz_when_PRF_l27_4_1 = 1'b0;
  assign _zz_when_PRF_l27_4 = {5'd0, _zz_when_PRF_l27_4_1};
  assign _zz_io_read_0_0_data_1 = io_read_0_0_idx;
  assign _zz_io_read_0_1_data_1 = io_read_0_1_idx;
  assign _zz_io_read_1_0_data_1 = io_read_1_0_idx;
  assign _zz_io_read_1_1_data_1 = io_read_1_1_idx;
  assign _zz_io_read_2_0_data_1 = io_read_2_0_idx;
  assign _zz_io_read_2_1_data_1 = io_read_2_1_idx;
  assign _zz_io_read_3_0_data_1 = io_read_3_0_idx;
  assign _zz_io_read_3_1_data_1 = io_read_3_1_idx;
  assign _zz_io_read_4_0_data_1 = io_read_4_0_idx;
  assign _zz_io_read_4_1_data_1 = io_read_4_1_idx;
  always @(*) begin
    case(_zz_io_read_0_0_data_1)
      6'b000000 : _zz_io_read_0_0_data = regFile_0;
      6'b000001 : _zz_io_read_0_0_data = regFile_1;
      6'b000010 : _zz_io_read_0_0_data = regFile_2;
      6'b000011 : _zz_io_read_0_0_data = regFile_3;
      6'b000100 : _zz_io_read_0_0_data = regFile_4;
      6'b000101 : _zz_io_read_0_0_data = regFile_5;
      6'b000110 : _zz_io_read_0_0_data = regFile_6;
      6'b000111 : _zz_io_read_0_0_data = regFile_7;
      6'b001000 : _zz_io_read_0_0_data = regFile_8;
      6'b001001 : _zz_io_read_0_0_data = regFile_9;
      6'b001010 : _zz_io_read_0_0_data = regFile_10;
      6'b001011 : _zz_io_read_0_0_data = regFile_11;
      6'b001100 : _zz_io_read_0_0_data = regFile_12;
      6'b001101 : _zz_io_read_0_0_data = regFile_13;
      6'b001110 : _zz_io_read_0_0_data = regFile_14;
      6'b001111 : _zz_io_read_0_0_data = regFile_15;
      6'b010000 : _zz_io_read_0_0_data = regFile_16;
      6'b010001 : _zz_io_read_0_0_data = regFile_17;
      6'b010010 : _zz_io_read_0_0_data = regFile_18;
      6'b010011 : _zz_io_read_0_0_data = regFile_19;
      6'b010100 : _zz_io_read_0_0_data = regFile_20;
      6'b010101 : _zz_io_read_0_0_data = regFile_21;
      6'b010110 : _zz_io_read_0_0_data = regFile_22;
      6'b010111 : _zz_io_read_0_0_data = regFile_23;
      6'b011000 : _zz_io_read_0_0_data = regFile_24;
      6'b011001 : _zz_io_read_0_0_data = regFile_25;
      6'b011010 : _zz_io_read_0_0_data = regFile_26;
      6'b011011 : _zz_io_read_0_0_data = regFile_27;
      6'b011100 : _zz_io_read_0_0_data = regFile_28;
      6'b011101 : _zz_io_read_0_0_data = regFile_29;
      6'b011110 : _zz_io_read_0_0_data = regFile_30;
      6'b011111 : _zz_io_read_0_0_data = regFile_31;
      6'b100000 : _zz_io_read_0_0_data = regFile_32;
      6'b100001 : _zz_io_read_0_0_data = regFile_33;
      6'b100010 : _zz_io_read_0_0_data = regFile_34;
      6'b100011 : _zz_io_read_0_0_data = regFile_35;
      6'b100100 : _zz_io_read_0_0_data = regFile_36;
      6'b100101 : _zz_io_read_0_0_data = regFile_37;
      6'b100110 : _zz_io_read_0_0_data = regFile_38;
      6'b100111 : _zz_io_read_0_0_data = regFile_39;
      6'b101000 : _zz_io_read_0_0_data = regFile_40;
      6'b101001 : _zz_io_read_0_0_data = regFile_41;
      6'b101010 : _zz_io_read_0_0_data = regFile_42;
      6'b101011 : _zz_io_read_0_0_data = regFile_43;
      6'b101100 : _zz_io_read_0_0_data = regFile_44;
      6'b101101 : _zz_io_read_0_0_data = regFile_45;
      6'b101110 : _zz_io_read_0_0_data = regFile_46;
      6'b101111 : _zz_io_read_0_0_data = regFile_47;
      6'b110000 : _zz_io_read_0_0_data = regFile_48;
      6'b110001 : _zz_io_read_0_0_data = regFile_49;
      6'b110010 : _zz_io_read_0_0_data = regFile_50;
      6'b110011 : _zz_io_read_0_0_data = regFile_51;
      6'b110100 : _zz_io_read_0_0_data = regFile_52;
      6'b110101 : _zz_io_read_0_0_data = regFile_53;
      6'b110110 : _zz_io_read_0_0_data = regFile_54;
      6'b110111 : _zz_io_read_0_0_data = regFile_55;
      6'b111000 : _zz_io_read_0_0_data = regFile_56;
      6'b111001 : _zz_io_read_0_0_data = regFile_57;
      6'b111010 : _zz_io_read_0_0_data = regFile_58;
      6'b111011 : _zz_io_read_0_0_data = regFile_59;
      6'b111100 : _zz_io_read_0_0_data = regFile_60;
      6'b111101 : _zz_io_read_0_0_data = regFile_61;
      6'b111110 : _zz_io_read_0_0_data = regFile_62;
      default : _zz_io_read_0_0_data = regFile_63;
    endcase
  end

  always @(*) begin
    case(_zz_io_read_0_1_data_1)
      6'b000000 : _zz_io_read_0_1_data = regFile_0;
      6'b000001 : _zz_io_read_0_1_data = regFile_1;
      6'b000010 : _zz_io_read_0_1_data = regFile_2;
      6'b000011 : _zz_io_read_0_1_data = regFile_3;
      6'b000100 : _zz_io_read_0_1_data = regFile_4;
      6'b000101 : _zz_io_read_0_1_data = regFile_5;
      6'b000110 : _zz_io_read_0_1_data = regFile_6;
      6'b000111 : _zz_io_read_0_1_data = regFile_7;
      6'b001000 : _zz_io_read_0_1_data = regFile_8;
      6'b001001 : _zz_io_read_0_1_data = regFile_9;
      6'b001010 : _zz_io_read_0_1_data = regFile_10;
      6'b001011 : _zz_io_read_0_1_data = regFile_11;
      6'b001100 : _zz_io_read_0_1_data = regFile_12;
      6'b001101 : _zz_io_read_0_1_data = regFile_13;
      6'b001110 : _zz_io_read_0_1_data = regFile_14;
      6'b001111 : _zz_io_read_0_1_data = regFile_15;
      6'b010000 : _zz_io_read_0_1_data = regFile_16;
      6'b010001 : _zz_io_read_0_1_data = regFile_17;
      6'b010010 : _zz_io_read_0_1_data = regFile_18;
      6'b010011 : _zz_io_read_0_1_data = regFile_19;
      6'b010100 : _zz_io_read_0_1_data = regFile_20;
      6'b010101 : _zz_io_read_0_1_data = regFile_21;
      6'b010110 : _zz_io_read_0_1_data = regFile_22;
      6'b010111 : _zz_io_read_0_1_data = regFile_23;
      6'b011000 : _zz_io_read_0_1_data = regFile_24;
      6'b011001 : _zz_io_read_0_1_data = regFile_25;
      6'b011010 : _zz_io_read_0_1_data = regFile_26;
      6'b011011 : _zz_io_read_0_1_data = regFile_27;
      6'b011100 : _zz_io_read_0_1_data = regFile_28;
      6'b011101 : _zz_io_read_0_1_data = regFile_29;
      6'b011110 : _zz_io_read_0_1_data = regFile_30;
      6'b011111 : _zz_io_read_0_1_data = regFile_31;
      6'b100000 : _zz_io_read_0_1_data = regFile_32;
      6'b100001 : _zz_io_read_0_1_data = regFile_33;
      6'b100010 : _zz_io_read_0_1_data = regFile_34;
      6'b100011 : _zz_io_read_0_1_data = regFile_35;
      6'b100100 : _zz_io_read_0_1_data = regFile_36;
      6'b100101 : _zz_io_read_0_1_data = regFile_37;
      6'b100110 : _zz_io_read_0_1_data = regFile_38;
      6'b100111 : _zz_io_read_0_1_data = regFile_39;
      6'b101000 : _zz_io_read_0_1_data = regFile_40;
      6'b101001 : _zz_io_read_0_1_data = regFile_41;
      6'b101010 : _zz_io_read_0_1_data = regFile_42;
      6'b101011 : _zz_io_read_0_1_data = regFile_43;
      6'b101100 : _zz_io_read_0_1_data = regFile_44;
      6'b101101 : _zz_io_read_0_1_data = regFile_45;
      6'b101110 : _zz_io_read_0_1_data = regFile_46;
      6'b101111 : _zz_io_read_0_1_data = regFile_47;
      6'b110000 : _zz_io_read_0_1_data = regFile_48;
      6'b110001 : _zz_io_read_0_1_data = regFile_49;
      6'b110010 : _zz_io_read_0_1_data = regFile_50;
      6'b110011 : _zz_io_read_0_1_data = regFile_51;
      6'b110100 : _zz_io_read_0_1_data = regFile_52;
      6'b110101 : _zz_io_read_0_1_data = regFile_53;
      6'b110110 : _zz_io_read_0_1_data = regFile_54;
      6'b110111 : _zz_io_read_0_1_data = regFile_55;
      6'b111000 : _zz_io_read_0_1_data = regFile_56;
      6'b111001 : _zz_io_read_0_1_data = regFile_57;
      6'b111010 : _zz_io_read_0_1_data = regFile_58;
      6'b111011 : _zz_io_read_0_1_data = regFile_59;
      6'b111100 : _zz_io_read_0_1_data = regFile_60;
      6'b111101 : _zz_io_read_0_1_data = regFile_61;
      6'b111110 : _zz_io_read_0_1_data = regFile_62;
      default : _zz_io_read_0_1_data = regFile_63;
    endcase
  end

  always @(*) begin
    case(_zz_io_read_1_0_data_1)
      6'b000000 : _zz_io_read_1_0_data = regFile_0;
      6'b000001 : _zz_io_read_1_0_data = regFile_1;
      6'b000010 : _zz_io_read_1_0_data = regFile_2;
      6'b000011 : _zz_io_read_1_0_data = regFile_3;
      6'b000100 : _zz_io_read_1_0_data = regFile_4;
      6'b000101 : _zz_io_read_1_0_data = regFile_5;
      6'b000110 : _zz_io_read_1_0_data = regFile_6;
      6'b000111 : _zz_io_read_1_0_data = regFile_7;
      6'b001000 : _zz_io_read_1_0_data = regFile_8;
      6'b001001 : _zz_io_read_1_0_data = regFile_9;
      6'b001010 : _zz_io_read_1_0_data = regFile_10;
      6'b001011 : _zz_io_read_1_0_data = regFile_11;
      6'b001100 : _zz_io_read_1_0_data = regFile_12;
      6'b001101 : _zz_io_read_1_0_data = regFile_13;
      6'b001110 : _zz_io_read_1_0_data = regFile_14;
      6'b001111 : _zz_io_read_1_0_data = regFile_15;
      6'b010000 : _zz_io_read_1_0_data = regFile_16;
      6'b010001 : _zz_io_read_1_0_data = regFile_17;
      6'b010010 : _zz_io_read_1_0_data = regFile_18;
      6'b010011 : _zz_io_read_1_0_data = regFile_19;
      6'b010100 : _zz_io_read_1_0_data = regFile_20;
      6'b010101 : _zz_io_read_1_0_data = regFile_21;
      6'b010110 : _zz_io_read_1_0_data = regFile_22;
      6'b010111 : _zz_io_read_1_0_data = regFile_23;
      6'b011000 : _zz_io_read_1_0_data = regFile_24;
      6'b011001 : _zz_io_read_1_0_data = regFile_25;
      6'b011010 : _zz_io_read_1_0_data = regFile_26;
      6'b011011 : _zz_io_read_1_0_data = regFile_27;
      6'b011100 : _zz_io_read_1_0_data = regFile_28;
      6'b011101 : _zz_io_read_1_0_data = regFile_29;
      6'b011110 : _zz_io_read_1_0_data = regFile_30;
      6'b011111 : _zz_io_read_1_0_data = regFile_31;
      6'b100000 : _zz_io_read_1_0_data = regFile_32;
      6'b100001 : _zz_io_read_1_0_data = regFile_33;
      6'b100010 : _zz_io_read_1_0_data = regFile_34;
      6'b100011 : _zz_io_read_1_0_data = regFile_35;
      6'b100100 : _zz_io_read_1_0_data = regFile_36;
      6'b100101 : _zz_io_read_1_0_data = regFile_37;
      6'b100110 : _zz_io_read_1_0_data = regFile_38;
      6'b100111 : _zz_io_read_1_0_data = regFile_39;
      6'b101000 : _zz_io_read_1_0_data = regFile_40;
      6'b101001 : _zz_io_read_1_0_data = regFile_41;
      6'b101010 : _zz_io_read_1_0_data = regFile_42;
      6'b101011 : _zz_io_read_1_0_data = regFile_43;
      6'b101100 : _zz_io_read_1_0_data = regFile_44;
      6'b101101 : _zz_io_read_1_0_data = regFile_45;
      6'b101110 : _zz_io_read_1_0_data = regFile_46;
      6'b101111 : _zz_io_read_1_0_data = regFile_47;
      6'b110000 : _zz_io_read_1_0_data = regFile_48;
      6'b110001 : _zz_io_read_1_0_data = regFile_49;
      6'b110010 : _zz_io_read_1_0_data = regFile_50;
      6'b110011 : _zz_io_read_1_0_data = regFile_51;
      6'b110100 : _zz_io_read_1_0_data = regFile_52;
      6'b110101 : _zz_io_read_1_0_data = regFile_53;
      6'b110110 : _zz_io_read_1_0_data = regFile_54;
      6'b110111 : _zz_io_read_1_0_data = regFile_55;
      6'b111000 : _zz_io_read_1_0_data = regFile_56;
      6'b111001 : _zz_io_read_1_0_data = regFile_57;
      6'b111010 : _zz_io_read_1_0_data = regFile_58;
      6'b111011 : _zz_io_read_1_0_data = regFile_59;
      6'b111100 : _zz_io_read_1_0_data = regFile_60;
      6'b111101 : _zz_io_read_1_0_data = regFile_61;
      6'b111110 : _zz_io_read_1_0_data = regFile_62;
      default : _zz_io_read_1_0_data = regFile_63;
    endcase
  end

  always @(*) begin
    case(_zz_io_read_1_1_data_1)
      6'b000000 : _zz_io_read_1_1_data = regFile_0;
      6'b000001 : _zz_io_read_1_1_data = regFile_1;
      6'b000010 : _zz_io_read_1_1_data = regFile_2;
      6'b000011 : _zz_io_read_1_1_data = regFile_3;
      6'b000100 : _zz_io_read_1_1_data = regFile_4;
      6'b000101 : _zz_io_read_1_1_data = regFile_5;
      6'b000110 : _zz_io_read_1_1_data = regFile_6;
      6'b000111 : _zz_io_read_1_1_data = regFile_7;
      6'b001000 : _zz_io_read_1_1_data = regFile_8;
      6'b001001 : _zz_io_read_1_1_data = regFile_9;
      6'b001010 : _zz_io_read_1_1_data = regFile_10;
      6'b001011 : _zz_io_read_1_1_data = regFile_11;
      6'b001100 : _zz_io_read_1_1_data = regFile_12;
      6'b001101 : _zz_io_read_1_1_data = regFile_13;
      6'b001110 : _zz_io_read_1_1_data = regFile_14;
      6'b001111 : _zz_io_read_1_1_data = regFile_15;
      6'b010000 : _zz_io_read_1_1_data = regFile_16;
      6'b010001 : _zz_io_read_1_1_data = regFile_17;
      6'b010010 : _zz_io_read_1_1_data = regFile_18;
      6'b010011 : _zz_io_read_1_1_data = regFile_19;
      6'b010100 : _zz_io_read_1_1_data = regFile_20;
      6'b010101 : _zz_io_read_1_1_data = regFile_21;
      6'b010110 : _zz_io_read_1_1_data = regFile_22;
      6'b010111 : _zz_io_read_1_1_data = regFile_23;
      6'b011000 : _zz_io_read_1_1_data = regFile_24;
      6'b011001 : _zz_io_read_1_1_data = regFile_25;
      6'b011010 : _zz_io_read_1_1_data = regFile_26;
      6'b011011 : _zz_io_read_1_1_data = regFile_27;
      6'b011100 : _zz_io_read_1_1_data = regFile_28;
      6'b011101 : _zz_io_read_1_1_data = regFile_29;
      6'b011110 : _zz_io_read_1_1_data = regFile_30;
      6'b011111 : _zz_io_read_1_1_data = regFile_31;
      6'b100000 : _zz_io_read_1_1_data = regFile_32;
      6'b100001 : _zz_io_read_1_1_data = regFile_33;
      6'b100010 : _zz_io_read_1_1_data = regFile_34;
      6'b100011 : _zz_io_read_1_1_data = regFile_35;
      6'b100100 : _zz_io_read_1_1_data = regFile_36;
      6'b100101 : _zz_io_read_1_1_data = regFile_37;
      6'b100110 : _zz_io_read_1_1_data = regFile_38;
      6'b100111 : _zz_io_read_1_1_data = regFile_39;
      6'b101000 : _zz_io_read_1_1_data = regFile_40;
      6'b101001 : _zz_io_read_1_1_data = regFile_41;
      6'b101010 : _zz_io_read_1_1_data = regFile_42;
      6'b101011 : _zz_io_read_1_1_data = regFile_43;
      6'b101100 : _zz_io_read_1_1_data = regFile_44;
      6'b101101 : _zz_io_read_1_1_data = regFile_45;
      6'b101110 : _zz_io_read_1_1_data = regFile_46;
      6'b101111 : _zz_io_read_1_1_data = regFile_47;
      6'b110000 : _zz_io_read_1_1_data = regFile_48;
      6'b110001 : _zz_io_read_1_1_data = regFile_49;
      6'b110010 : _zz_io_read_1_1_data = regFile_50;
      6'b110011 : _zz_io_read_1_1_data = regFile_51;
      6'b110100 : _zz_io_read_1_1_data = regFile_52;
      6'b110101 : _zz_io_read_1_1_data = regFile_53;
      6'b110110 : _zz_io_read_1_1_data = regFile_54;
      6'b110111 : _zz_io_read_1_1_data = regFile_55;
      6'b111000 : _zz_io_read_1_1_data = regFile_56;
      6'b111001 : _zz_io_read_1_1_data = regFile_57;
      6'b111010 : _zz_io_read_1_1_data = regFile_58;
      6'b111011 : _zz_io_read_1_1_data = regFile_59;
      6'b111100 : _zz_io_read_1_1_data = regFile_60;
      6'b111101 : _zz_io_read_1_1_data = regFile_61;
      6'b111110 : _zz_io_read_1_1_data = regFile_62;
      default : _zz_io_read_1_1_data = regFile_63;
    endcase
  end

  always @(*) begin
    case(_zz_io_read_2_0_data_1)
      6'b000000 : _zz_io_read_2_0_data = regFile_0;
      6'b000001 : _zz_io_read_2_0_data = regFile_1;
      6'b000010 : _zz_io_read_2_0_data = regFile_2;
      6'b000011 : _zz_io_read_2_0_data = regFile_3;
      6'b000100 : _zz_io_read_2_0_data = regFile_4;
      6'b000101 : _zz_io_read_2_0_data = regFile_5;
      6'b000110 : _zz_io_read_2_0_data = regFile_6;
      6'b000111 : _zz_io_read_2_0_data = regFile_7;
      6'b001000 : _zz_io_read_2_0_data = regFile_8;
      6'b001001 : _zz_io_read_2_0_data = regFile_9;
      6'b001010 : _zz_io_read_2_0_data = regFile_10;
      6'b001011 : _zz_io_read_2_0_data = regFile_11;
      6'b001100 : _zz_io_read_2_0_data = regFile_12;
      6'b001101 : _zz_io_read_2_0_data = regFile_13;
      6'b001110 : _zz_io_read_2_0_data = regFile_14;
      6'b001111 : _zz_io_read_2_0_data = regFile_15;
      6'b010000 : _zz_io_read_2_0_data = regFile_16;
      6'b010001 : _zz_io_read_2_0_data = regFile_17;
      6'b010010 : _zz_io_read_2_0_data = regFile_18;
      6'b010011 : _zz_io_read_2_0_data = regFile_19;
      6'b010100 : _zz_io_read_2_0_data = regFile_20;
      6'b010101 : _zz_io_read_2_0_data = regFile_21;
      6'b010110 : _zz_io_read_2_0_data = regFile_22;
      6'b010111 : _zz_io_read_2_0_data = regFile_23;
      6'b011000 : _zz_io_read_2_0_data = regFile_24;
      6'b011001 : _zz_io_read_2_0_data = regFile_25;
      6'b011010 : _zz_io_read_2_0_data = regFile_26;
      6'b011011 : _zz_io_read_2_0_data = regFile_27;
      6'b011100 : _zz_io_read_2_0_data = regFile_28;
      6'b011101 : _zz_io_read_2_0_data = regFile_29;
      6'b011110 : _zz_io_read_2_0_data = regFile_30;
      6'b011111 : _zz_io_read_2_0_data = regFile_31;
      6'b100000 : _zz_io_read_2_0_data = regFile_32;
      6'b100001 : _zz_io_read_2_0_data = regFile_33;
      6'b100010 : _zz_io_read_2_0_data = regFile_34;
      6'b100011 : _zz_io_read_2_0_data = regFile_35;
      6'b100100 : _zz_io_read_2_0_data = regFile_36;
      6'b100101 : _zz_io_read_2_0_data = regFile_37;
      6'b100110 : _zz_io_read_2_0_data = regFile_38;
      6'b100111 : _zz_io_read_2_0_data = regFile_39;
      6'b101000 : _zz_io_read_2_0_data = regFile_40;
      6'b101001 : _zz_io_read_2_0_data = regFile_41;
      6'b101010 : _zz_io_read_2_0_data = regFile_42;
      6'b101011 : _zz_io_read_2_0_data = regFile_43;
      6'b101100 : _zz_io_read_2_0_data = regFile_44;
      6'b101101 : _zz_io_read_2_0_data = regFile_45;
      6'b101110 : _zz_io_read_2_0_data = regFile_46;
      6'b101111 : _zz_io_read_2_0_data = regFile_47;
      6'b110000 : _zz_io_read_2_0_data = regFile_48;
      6'b110001 : _zz_io_read_2_0_data = regFile_49;
      6'b110010 : _zz_io_read_2_0_data = regFile_50;
      6'b110011 : _zz_io_read_2_0_data = regFile_51;
      6'b110100 : _zz_io_read_2_0_data = regFile_52;
      6'b110101 : _zz_io_read_2_0_data = regFile_53;
      6'b110110 : _zz_io_read_2_0_data = regFile_54;
      6'b110111 : _zz_io_read_2_0_data = regFile_55;
      6'b111000 : _zz_io_read_2_0_data = regFile_56;
      6'b111001 : _zz_io_read_2_0_data = regFile_57;
      6'b111010 : _zz_io_read_2_0_data = regFile_58;
      6'b111011 : _zz_io_read_2_0_data = regFile_59;
      6'b111100 : _zz_io_read_2_0_data = regFile_60;
      6'b111101 : _zz_io_read_2_0_data = regFile_61;
      6'b111110 : _zz_io_read_2_0_data = regFile_62;
      default : _zz_io_read_2_0_data = regFile_63;
    endcase
  end

  always @(*) begin
    case(_zz_io_read_2_1_data_1)
      6'b000000 : _zz_io_read_2_1_data = regFile_0;
      6'b000001 : _zz_io_read_2_1_data = regFile_1;
      6'b000010 : _zz_io_read_2_1_data = regFile_2;
      6'b000011 : _zz_io_read_2_1_data = regFile_3;
      6'b000100 : _zz_io_read_2_1_data = regFile_4;
      6'b000101 : _zz_io_read_2_1_data = regFile_5;
      6'b000110 : _zz_io_read_2_1_data = regFile_6;
      6'b000111 : _zz_io_read_2_1_data = regFile_7;
      6'b001000 : _zz_io_read_2_1_data = regFile_8;
      6'b001001 : _zz_io_read_2_1_data = regFile_9;
      6'b001010 : _zz_io_read_2_1_data = regFile_10;
      6'b001011 : _zz_io_read_2_1_data = regFile_11;
      6'b001100 : _zz_io_read_2_1_data = regFile_12;
      6'b001101 : _zz_io_read_2_1_data = regFile_13;
      6'b001110 : _zz_io_read_2_1_data = regFile_14;
      6'b001111 : _zz_io_read_2_1_data = regFile_15;
      6'b010000 : _zz_io_read_2_1_data = regFile_16;
      6'b010001 : _zz_io_read_2_1_data = regFile_17;
      6'b010010 : _zz_io_read_2_1_data = regFile_18;
      6'b010011 : _zz_io_read_2_1_data = regFile_19;
      6'b010100 : _zz_io_read_2_1_data = regFile_20;
      6'b010101 : _zz_io_read_2_1_data = regFile_21;
      6'b010110 : _zz_io_read_2_1_data = regFile_22;
      6'b010111 : _zz_io_read_2_1_data = regFile_23;
      6'b011000 : _zz_io_read_2_1_data = regFile_24;
      6'b011001 : _zz_io_read_2_1_data = regFile_25;
      6'b011010 : _zz_io_read_2_1_data = regFile_26;
      6'b011011 : _zz_io_read_2_1_data = regFile_27;
      6'b011100 : _zz_io_read_2_1_data = regFile_28;
      6'b011101 : _zz_io_read_2_1_data = regFile_29;
      6'b011110 : _zz_io_read_2_1_data = regFile_30;
      6'b011111 : _zz_io_read_2_1_data = regFile_31;
      6'b100000 : _zz_io_read_2_1_data = regFile_32;
      6'b100001 : _zz_io_read_2_1_data = regFile_33;
      6'b100010 : _zz_io_read_2_1_data = regFile_34;
      6'b100011 : _zz_io_read_2_1_data = regFile_35;
      6'b100100 : _zz_io_read_2_1_data = regFile_36;
      6'b100101 : _zz_io_read_2_1_data = regFile_37;
      6'b100110 : _zz_io_read_2_1_data = regFile_38;
      6'b100111 : _zz_io_read_2_1_data = regFile_39;
      6'b101000 : _zz_io_read_2_1_data = regFile_40;
      6'b101001 : _zz_io_read_2_1_data = regFile_41;
      6'b101010 : _zz_io_read_2_1_data = regFile_42;
      6'b101011 : _zz_io_read_2_1_data = regFile_43;
      6'b101100 : _zz_io_read_2_1_data = regFile_44;
      6'b101101 : _zz_io_read_2_1_data = regFile_45;
      6'b101110 : _zz_io_read_2_1_data = regFile_46;
      6'b101111 : _zz_io_read_2_1_data = regFile_47;
      6'b110000 : _zz_io_read_2_1_data = regFile_48;
      6'b110001 : _zz_io_read_2_1_data = regFile_49;
      6'b110010 : _zz_io_read_2_1_data = regFile_50;
      6'b110011 : _zz_io_read_2_1_data = regFile_51;
      6'b110100 : _zz_io_read_2_1_data = regFile_52;
      6'b110101 : _zz_io_read_2_1_data = regFile_53;
      6'b110110 : _zz_io_read_2_1_data = regFile_54;
      6'b110111 : _zz_io_read_2_1_data = regFile_55;
      6'b111000 : _zz_io_read_2_1_data = regFile_56;
      6'b111001 : _zz_io_read_2_1_data = regFile_57;
      6'b111010 : _zz_io_read_2_1_data = regFile_58;
      6'b111011 : _zz_io_read_2_1_data = regFile_59;
      6'b111100 : _zz_io_read_2_1_data = regFile_60;
      6'b111101 : _zz_io_read_2_1_data = regFile_61;
      6'b111110 : _zz_io_read_2_1_data = regFile_62;
      default : _zz_io_read_2_1_data = regFile_63;
    endcase
  end

  always @(*) begin
    case(_zz_io_read_3_0_data_1)
      6'b000000 : _zz_io_read_3_0_data = regFile_0;
      6'b000001 : _zz_io_read_3_0_data = regFile_1;
      6'b000010 : _zz_io_read_3_0_data = regFile_2;
      6'b000011 : _zz_io_read_3_0_data = regFile_3;
      6'b000100 : _zz_io_read_3_0_data = regFile_4;
      6'b000101 : _zz_io_read_3_0_data = regFile_5;
      6'b000110 : _zz_io_read_3_0_data = regFile_6;
      6'b000111 : _zz_io_read_3_0_data = regFile_7;
      6'b001000 : _zz_io_read_3_0_data = regFile_8;
      6'b001001 : _zz_io_read_3_0_data = regFile_9;
      6'b001010 : _zz_io_read_3_0_data = regFile_10;
      6'b001011 : _zz_io_read_3_0_data = regFile_11;
      6'b001100 : _zz_io_read_3_0_data = regFile_12;
      6'b001101 : _zz_io_read_3_0_data = regFile_13;
      6'b001110 : _zz_io_read_3_0_data = regFile_14;
      6'b001111 : _zz_io_read_3_0_data = regFile_15;
      6'b010000 : _zz_io_read_3_0_data = regFile_16;
      6'b010001 : _zz_io_read_3_0_data = regFile_17;
      6'b010010 : _zz_io_read_3_0_data = regFile_18;
      6'b010011 : _zz_io_read_3_0_data = regFile_19;
      6'b010100 : _zz_io_read_3_0_data = regFile_20;
      6'b010101 : _zz_io_read_3_0_data = regFile_21;
      6'b010110 : _zz_io_read_3_0_data = regFile_22;
      6'b010111 : _zz_io_read_3_0_data = regFile_23;
      6'b011000 : _zz_io_read_3_0_data = regFile_24;
      6'b011001 : _zz_io_read_3_0_data = regFile_25;
      6'b011010 : _zz_io_read_3_0_data = regFile_26;
      6'b011011 : _zz_io_read_3_0_data = regFile_27;
      6'b011100 : _zz_io_read_3_0_data = regFile_28;
      6'b011101 : _zz_io_read_3_0_data = regFile_29;
      6'b011110 : _zz_io_read_3_0_data = regFile_30;
      6'b011111 : _zz_io_read_3_0_data = regFile_31;
      6'b100000 : _zz_io_read_3_0_data = regFile_32;
      6'b100001 : _zz_io_read_3_0_data = regFile_33;
      6'b100010 : _zz_io_read_3_0_data = regFile_34;
      6'b100011 : _zz_io_read_3_0_data = regFile_35;
      6'b100100 : _zz_io_read_3_0_data = regFile_36;
      6'b100101 : _zz_io_read_3_0_data = regFile_37;
      6'b100110 : _zz_io_read_3_0_data = regFile_38;
      6'b100111 : _zz_io_read_3_0_data = regFile_39;
      6'b101000 : _zz_io_read_3_0_data = regFile_40;
      6'b101001 : _zz_io_read_3_0_data = regFile_41;
      6'b101010 : _zz_io_read_3_0_data = regFile_42;
      6'b101011 : _zz_io_read_3_0_data = regFile_43;
      6'b101100 : _zz_io_read_3_0_data = regFile_44;
      6'b101101 : _zz_io_read_3_0_data = regFile_45;
      6'b101110 : _zz_io_read_3_0_data = regFile_46;
      6'b101111 : _zz_io_read_3_0_data = regFile_47;
      6'b110000 : _zz_io_read_3_0_data = regFile_48;
      6'b110001 : _zz_io_read_3_0_data = regFile_49;
      6'b110010 : _zz_io_read_3_0_data = regFile_50;
      6'b110011 : _zz_io_read_3_0_data = regFile_51;
      6'b110100 : _zz_io_read_3_0_data = regFile_52;
      6'b110101 : _zz_io_read_3_0_data = regFile_53;
      6'b110110 : _zz_io_read_3_0_data = regFile_54;
      6'b110111 : _zz_io_read_3_0_data = regFile_55;
      6'b111000 : _zz_io_read_3_0_data = regFile_56;
      6'b111001 : _zz_io_read_3_0_data = regFile_57;
      6'b111010 : _zz_io_read_3_0_data = regFile_58;
      6'b111011 : _zz_io_read_3_0_data = regFile_59;
      6'b111100 : _zz_io_read_3_0_data = regFile_60;
      6'b111101 : _zz_io_read_3_0_data = regFile_61;
      6'b111110 : _zz_io_read_3_0_data = regFile_62;
      default : _zz_io_read_3_0_data = regFile_63;
    endcase
  end

  always @(*) begin
    case(_zz_io_read_3_1_data_1)
      6'b000000 : _zz_io_read_3_1_data = regFile_0;
      6'b000001 : _zz_io_read_3_1_data = regFile_1;
      6'b000010 : _zz_io_read_3_1_data = regFile_2;
      6'b000011 : _zz_io_read_3_1_data = regFile_3;
      6'b000100 : _zz_io_read_3_1_data = regFile_4;
      6'b000101 : _zz_io_read_3_1_data = regFile_5;
      6'b000110 : _zz_io_read_3_1_data = regFile_6;
      6'b000111 : _zz_io_read_3_1_data = regFile_7;
      6'b001000 : _zz_io_read_3_1_data = regFile_8;
      6'b001001 : _zz_io_read_3_1_data = regFile_9;
      6'b001010 : _zz_io_read_3_1_data = regFile_10;
      6'b001011 : _zz_io_read_3_1_data = regFile_11;
      6'b001100 : _zz_io_read_3_1_data = regFile_12;
      6'b001101 : _zz_io_read_3_1_data = regFile_13;
      6'b001110 : _zz_io_read_3_1_data = regFile_14;
      6'b001111 : _zz_io_read_3_1_data = regFile_15;
      6'b010000 : _zz_io_read_3_1_data = regFile_16;
      6'b010001 : _zz_io_read_3_1_data = regFile_17;
      6'b010010 : _zz_io_read_3_1_data = regFile_18;
      6'b010011 : _zz_io_read_3_1_data = regFile_19;
      6'b010100 : _zz_io_read_3_1_data = regFile_20;
      6'b010101 : _zz_io_read_3_1_data = regFile_21;
      6'b010110 : _zz_io_read_3_1_data = regFile_22;
      6'b010111 : _zz_io_read_3_1_data = regFile_23;
      6'b011000 : _zz_io_read_3_1_data = regFile_24;
      6'b011001 : _zz_io_read_3_1_data = regFile_25;
      6'b011010 : _zz_io_read_3_1_data = regFile_26;
      6'b011011 : _zz_io_read_3_1_data = regFile_27;
      6'b011100 : _zz_io_read_3_1_data = regFile_28;
      6'b011101 : _zz_io_read_3_1_data = regFile_29;
      6'b011110 : _zz_io_read_3_1_data = regFile_30;
      6'b011111 : _zz_io_read_3_1_data = regFile_31;
      6'b100000 : _zz_io_read_3_1_data = regFile_32;
      6'b100001 : _zz_io_read_3_1_data = regFile_33;
      6'b100010 : _zz_io_read_3_1_data = regFile_34;
      6'b100011 : _zz_io_read_3_1_data = regFile_35;
      6'b100100 : _zz_io_read_3_1_data = regFile_36;
      6'b100101 : _zz_io_read_3_1_data = regFile_37;
      6'b100110 : _zz_io_read_3_1_data = regFile_38;
      6'b100111 : _zz_io_read_3_1_data = regFile_39;
      6'b101000 : _zz_io_read_3_1_data = regFile_40;
      6'b101001 : _zz_io_read_3_1_data = regFile_41;
      6'b101010 : _zz_io_read_3_1_data = regFile_42;
      6'b101011 : _zz_io_read_3_1_data = regFile_43;
      6'b101100 : _zz_io_read_3_1_data = regFile_44;
      6'b101101 : _zz_io_read_3_1_data = regFile_45;
      6'b101110 : _zz_io_read_3_1_data = regFile_46;
      6'b101111 : _zz_io_read_3_1_data = regFile_47;
      6'b110000 : _zz_io_read_3_1_data = regFile_48;
      6'b110001 : _zz_io_read_3_1_data = regFile_49;
      6'b110010 : _zz_io_read_3_1_data = regFile_50;
      6'b110011 : _zz_io_read_3_1_data = regFile_51;
      6'b110100 : _zz_io_read_3_1_data = regFile_52;
      6'b110101 : _zz_io_read_3_1_data = regFile_53;
      6'b110110 : _zz_io_read_3_1_data = regFile_54;
      6'b110111 : _zz_io_read_3_1_data = regFile_55;
      6'b111000 : _zz_io_read_3_1_data = regFile_56;
      6'b111001 : _zz_io_read_3_1_data = regFile_57;
      6'b111010 : _zz_io_read_3_1_data = regFile_58;
      6'b111011 : _zz_io_read_3_1_data = regFile_59;
      6'b111100 : _zz_io_read_3_1_data = regFile_60;
      6'b111101 : _zz_io_read_3_1_data = regFile_61;
      6'b111110 : _zz_io_read_3_1_data = regFile_62;
      default : _zz_io_read_3_1_data = regFile_63;
    endcase
  end

  always @(*) begin
    case(_zz_io_read_4_0_data_1)
      6'b000000 : _zz_io_read_4_0_data = regFile_0;
      6'b000001 : _zz_io_read_4_0_data = regFile_1;
      6'b000010 : _zz_io_read_4_0_data = regFile_2;
      6'b000011 : _zz_io_read_4_0_data = regFile_3;
      6'b000100 : _zz_io_read_4_0_data = regFile_4;
      6'b000101 : _zz_io_read_4_0_data = regFile_5;
      6'b000110 : _zz_io_read_4_0_data = regFile_6;
      6'b000111 : _zz_io_read_4_0_data = regFile_7;
      6'b001000 : _zz_io_read_4_0_data = regFile_8;
      6'b001001 : _zz_io_read_4_0_data = regFile_9;
      6'b001010 : _zz_io_read_4_0_data = regFile_10;
      6'b001011 : _zz_io_read_4_0_data = regFile_11;
      6'b001100 : _zz_io_read_4_0_data = regFile_12;
      6'b001101 : _zz_io_read_4_0_data = regFile_13;
      6'b001110 : _zz_io_read_4_0_data = regFile_14;
      6'b001111 : _zz_io_read_4_0_data = regFile_15;
      6'b010000 : _zz_io_read_4_0_data = regFile_16;
      6'b010001 : _zz_io_read_4_0_data = regFile_17;
      6'b010010 : _zz_io_read_4_0_data = regFile_18;
      6'b010011 : _zz_io_read_4_0_data = regFile_19;
      6'b010100 : _zz_io_read_4_0_data = regFile_20;
      6'b010101 : _zz_io_read_4_0_data = regFile_21;
      6'b010110 : _zz_io_read_4_0_data = regFile_22;
      6'b010111 : _zz_io_read_4_0_data = regFile_23;
      6'b011000 : _zz_io_read_4_0_data = regFile_24;
      6'b011001 : _zz_io_read_4_0_data = regFile_25;
      6'b011010 : _zz_io_read_4_0_data = regFile_26;
      6'b011011 : _zz_io_read_4_0_data = regFile_27;
      6'b011100 : _zz_io_read_4_0_data = regFile_28;
      6'b011101 : _zz_io_read_4_0_data = regFile_29;
      6'b011110 : _zz_io_read_4_0_data = regFile_30;
      6'b011111 : _zz_io_read_4_0_data = regFile_31;
      6'b100000 : _zz_io_read_4_0_data = regFile_32;
      6'b100001 : _zz_io_read_4_0_data = regFile_33;
      6'b100010 : _zz_io_read_4_0_data = regFile_34;
      6'b100011 : _zz_io_read_4_0_data = regFile_35;
      6'b100100 : _zz_io_read_4_0_data = regFile_36;
      6'b100101 : _zz_io_read_4_0_data = regFile_37;
      6'b100110 : _zz_io_read_4_0_data = regFile_38;
      6'b100111 : _zz_io_read_4_0_data = regFile_39;
      6'b101000 : _zz_io_read_4_0_data = regFile_40;
      6'b101001 : _zz_io_read_4_0_data = regFile_41;
      6'b101010 : _zz_io_read_4_0_data = regFile_42;
      6'b101011 : _zz_io_read_4_0_data = regFile_43;
      6'b101100 : _zz_io_read_4_0_data = regFile_44;
      6'b101101 : _zz_io_read_4_0_data = regFile_45;
      6'b101110 : _zz_io_read_4_0_data = regFile_46;
      6'b101111 : _zz_io_read_4_0_data = regFile_47;
      6'b110000 : _zz_io_read_4_0_data = regFile_48;
      6'b110001 : _zz_io_read_4_0_data = regFile_49;
      6'b110010 : _zz_io_read_4_0_data = regFile_50;
      6'b110011 : _zz_io_read_4_0_data = regFile_51;
      6'b110100 : _zz_io_read_4_0_data = regFile_52;
      6'b110101 : _zz_io_read_4_0_data = regFile_53;
      6'b110110 : _zz_io_read_4_0_data = regFile_54;
      6'b110111 : _zz_io_read_4_0_data = regFile_55;
      6'b111000 : _zz_io_read_4_0_data = regFile_56;
      6'b111001 : _zz_io_read_4_0_data = regFile_57;
      6'b111010 : _zz_io_read_4_0_data = regFile_58;
      6'b111011 : _zz_io_read_4_0_data = regFile_59;
      6'b111100 : _zz_io_read_4_0_data = regFile_60;
      6'b111101 : _zz_io_read_4_0_data = regFile_61;
      6'b111110 : _zz_io_read_4_0_data = regFile_62;
      default : _zz_io_read_4_0_data = regFile_63;
    endcase
  end

  always @(*) begin
    case(_zz_io_read_4_1_data_1)
      6'b000000 : _zz_io_read_4_1_data = regFile_0;
      6'b000001 : _zz_io_read_4_1_data = regFile_1;
      6'b000010 : _zz_io_read_4_1_data = regFile_2;
      6'b000011 : _zz_io_read_4_1_data = regFile_3;
      6'b000100 : _zz_io_read_4_1_data = regFile_4;
      6'b000101 : _zz_io_read_4_1_data = regFile_5;
      6'b000110 : _zz_io_read_4_1_data = regFile_6;
      6'b000111 : _zz_io_read_4_1_data = regFile_7;
      6'b001000 : _zz_io_read_4_1_data = regFile_8;
      6'b001001 : _zz_io_read_4_1_data = regFile_9;
      6'b001010 : _zz_io_read_4_1_data = regFile_10;
      6'b001011 : _zz_io_read_4_1_data = regFile_11;
      6'b001100 : _zz_io_read_4_1_data = regFile_12;
      6'b001101 : _zz_io_read_4_1_data = regFile_13;
      6'b001110 : _zz_io_read_4_1_data = regFile_14;
      6'b001111 : _zz_io_read_4_1_data = regFile_15;
      6'b010000 : _zz_io_read_4_1_data = regFile_16;
      6'b010001 : _zz_io_read_4_1_data = regFile_17;
      6'b010010 : _zz_io_read_4_1_data = regFile_18;
      6'b010011 : _zz_io_read_4_1_data = regFile_19;
      6'b010100 : _zz_io_read_4_1_data = regFile_20;
      6'b010101 : _zz_io_read_4_1_data = regFile_21;
      6'b010110 : _zz_io_read_4_1_data = regFile_22;
      6'b010111 : _zz_io_read_4_1_data = regFile_23;
      6'b011000 : _zz_io_read_4_1_data = regFile_24;
      6'b011001 : _zz_io_read_4_1_data = regFile_25;
      6'b011010 : _zz_io_read_4_1_data = regFile_26;
      6'b011011 : _zz_io_read_4_1_data = regFile_27;
      6'b011100 : _zz_io_read_4_1_data = regFile_28;
      6'b011101 : _zz_io_read_4_1_data = regFile_29;
      6'b011110 : _zz_io_read_4_1_data = regFile_30;
      6'b011111 : _zz_io_read_4_1_data = regFile_31;
      6'b100000 : _zz_io_read_4_1_data = regFile_32;
      6'b100001 : _zz_io_read_4_1_data = regFile_33;
      6'b100010 : _zz_io_read_4_1_data = regFile_34;
      6'b100011 : _zz_io_read_4_1_data = regFile_35;
      6'b100100 : _zz_io_read_4_1_data = regFile_36;
      6'b100101 : _zz_io_read_4_1_data = regFile_37;
      6'b100110 : _zz_io_read_4_1_data = regFile_38;
      6'b100111 : _zz_io_read_4_1_data = regFile_39;
      6'b101000 : _zz_io_read_4_1_data = regFile_40;
      6'b101001 : _zz_io_read_4_1_data = regFile_41;
      6'b101010 : _zz_io_read_4_1_data = regFile_42;
      6'b101011 : _zz_io_read_4_1_data = regFile_43;
      6'b101100 : _zz_io_read_4_1_data = regFile_44;
      6'b101101 : _zz_io_read_4_1_data = regFile_45;
      6'b101110 : _zz_io_read_4_1_data = regFile_46;
      6'b101111 : _zz_io_read_4_1_data = regFile_47;
      6'b110000 : _zz_io_read_4_1_data = regFile_48;
      6'b110001 : _zz_io_read_4_1_data = regFile_49;
      6'b110010 : _zz_io_read_4_1_data = regFile_50;
      6'b110011 : _zz_io_read_4_1_data = regFile_51;
      6'b110100 : _zz_io_read_4_1_data = regFile_52;
      6'b110101 : _zz_io_read_4_1_data = regFile_53;
      6'b110110 : _zz_io_read_4_1_data = regFile_54;
      6'b110111 : _zz_io_read_4_1_data = regFile_55;
      6'b111000 : _zz_io_read_4_1_data = regFile_56;
      6'b111001 : _zz_io_read_4_1_data = regFile_57;
      6'b111010 : _zz_io_read_4_1_data = regFile_58;
      6'b111011 : _zz_io_read_4_1_data = regFile_59;
      6'b111100 : _zz_io_read_4_1_data = regFile_60;
      6'b111101 : _zz_io_read_4_1_data = regFile_61;
      6'b111110 : _zz_io_read_4_1_data = regFile_62;
      default : _zz_io_read_4_1_data = regFile_63;
    endcase
  end

  assign when_PRF_l19 = (io_read_0_0_idx != _zz_when_PRF_l19);
  always @(*) begin
    if(when_PRF_l19) begin
      io_read_0_0_data = _zz_io_read_0_0_data;
    end else begin
      io_read_0_0_data = {31'd0, _zz_io_read_0_0_data_2};
    end
  end

  assign when_PRF_l19_1 = (io_read_0_1_idx != _zz_when_PRF_l19_1_1);
  always @(*) begin
    if(when_PRF_l19_1) begin
      io_read_0_1_data = _zz_io_read_0_1_data;
    end else begin
      io_read_0_1_data = {31'd0, _zz_io_read_0_1_data_2};
    end
  end

  assign when_PRF_l19_2 = (io_read_1_0_idx != _zz_when_PRF_l19_2);
  always @(*) begin
    if(when_PRF_l19_2) begin
      io_read_1_0_data = _zz_io_read_1_0_data;
    end else begin
      io_read_1_0_data = {31'd0, _zz_io_read_1_0_data_2};
    end
  end

  assign when_PRF_l19_3 = (io_read_1_1_idx != _zz_when_PRF_l19_3);
  always @(*) begin
    if(when_PRF_l19_3) begin
      io_read_1_1_data = _zz_io_read_1_1_data;
    end else begin
      io_read_1_1_data = {31'd0, _zz_io_read_1_1_data_2};
    end
  end

  assign when_PRF_l19_4 = (io_read_2_0_idx != _zz_when_PRF_l19_4);
  always @(*) begin
    if(when_PRF_l19_4) begin
      io_read_2_0_data = _zz_io_read_2_0_data;
    end else begin
      io_read_2_0_data = {31'd0, _zz_io_read_2_0_data_2};
    end
  end

  assign when_PRF_l19_5 = (io_read_2_1_idx != _zz_when_PRF_l19_5);
  always @(*) begin
    if(when_PRF_l19_5) begin
      io_read_2_1_data = _zz_io_read_2_1_data;
    end else begin
      io_read_2_1_data = {31'd0, _zz_io_read_2_1_data_2};
    end
  end

  assign when_PRF_l19_6 = (io_read_3_0_idx != _zz_when_PRF_l19_6);
  always @(*) begin
    if(when_PRF_l19_6) begin
      io_read_3_0_data = _zz_io_read_3_0_data;
    end else begin
      io_read_3_0_data = {31'd0, _zz_io_read_3_0_data_2};
    end
  end

  assign when_PRF_l19_7 = (io_read_3_1_idx != _zz_when_PRF_l19_7);
  always @(*) begin
    if(when_PRF_l19_7) begin
      io_read_3_1_data = _zz_io_read_3_1_data;
    end else begin
      io_read_3_1_data = {31'd0, _zz_io_read_3_1_data_2};
    end
  end

  assign when_PRF_l19_8 = (io_read_4_0_idx != _zz_when_PRF_l19_8);
  always @(*) begin
    if(when_PRF_l19_8) begin
      io_read_4_0_data = _zz_io_read_4_0_data;
    end else begin
      io_read_4_0_data = {31'd0, _zz_io_read_4_0_data_2};
    end
  end

  assign when_PRF_l19_9 = (io_read_4_1_idx != _zz_when_PRF_l19_9);
  always @(*) begin
    if(when_PRF_l19_9) begin
      io_read_4_1_data = _zz_io_read_4_1_data;
    end else begin
      io_read_4_1_data = {31'd0, _zz_io_read_4_1_data_2};
    end
  end

  assign when_PRF_l27 = (io_write_0_idx != _zz_when_PRF_l27);
  assign _zz_1 = ({63'd0,1'b1} <<< io_write_0_idx);
  assign when_PRF_l27_1 = (io_write_1_idx != _zz_when_PRF_l27_1_1);
  assign _zz_2 = ({63'd0,1'b1} <<< io_write_1_idx);
  assign when_PRF_l27_2 = (io_write_2_idx != _zz_when_PRF_l27_2);
  assign _zz_3 = ({63'd0,1'b1} <<< io_write_2_idx);
  assign when_PRF_l27_3 = (io_write_3_idx != _zz_when_PRF_l27_3);
  assign _zz_4 = ({63'd0,1'b1} <<< io_write_3_idx);
  assign when_PRF_l27_4 = (io_write_4_idx != _zz_when_PRF_l27_4);
  assign _zz_5 = ({63'd0,1'b1} <<< io_write_4_idx);
  always @(posedge aclk) begin
    if(when_PRF_l27) begin
      if(_zz_1[0]) begin
        regFile_0 <= io_write_0_data;
      end
      if(_zz_1[1]) begin
        regFile_1 <= io_write_0_data;
      end
      if(_zz_1[2]) begin
        regFile_2 <= io_write_0_data;
      end
      if(_zz_1[3]) begin
        regFile_3 <= io_write_0_data;
      end
      if(_zz_1[4]) begin
        regFile_4 <= io_write_0_data;
      end
      if(_zz_1[5]) begin
        regFile_5 <= io_write_0_data;
      end
      if(_zz_1[6]) begin
        regFile_6 <= io_write_0_data;
      end
      if(_zz_1[7]) begin
        regFile_7 <= io_write_0_data;
      end
      if(_zz_1[8]) begin
        regFile_8 <= io_write_0_data;
      end
      if(_zz_1[9]) begin
        regFile_9 <= io_write_0_data;
      end
      if(_zz_1[10]) begin
        regFile_10 <= io_write_0_data;
      end
      if(_zz_1[11]) begin
        regFile_11 <= io_write_0_data;
      end
      if(_zz_1[12]) begin
        regFile_12 <= io_write_0_data;
      end
      if(_zz_1[13]) begin
        regFile_13 <= io_write_0_data;
      end
      if(_zz_1[14]) begin
        regFile_14 <= io_write_0_data;
      end
      if(_zz_1[15]) begin
        regFile_15 <= io_write_0_data;
      end
      if(_zz_1[16]) begin
        regFile_16 <= io_write_0_data;
      end
      if(_zz_1[17]) begin
        regFile_17 <= io_write_0_data;
      end
      if(_zz_1[18]) begin
        regFile_18 <= io_write_0_data;
      end
      if(_zz_1[19]) begin
        regFile_19 <= io_write_0_data;
      end
      if(_zz_1[20]) begin
        regFile_20 <= io_write_0_data;
      end
      if(_zz_1[21]) begin
        regFile_21 <= io_write_0_data;
      end
      if(_zz_1[22]) begin
        regFile_22 <= io_write_0_data;
      end
      if(_zz_1[23]) begin
        regFile_23 <= io_write_0_data;
      end
      if(_zz_1[24]) begin
        regFile_24 <= io_write_0_data;
      end
      if(_zz_1[25]) begin
        regFile_25 <= io_write_0_data;
      end
      if(_zz_1[26]) begin
        regFile_26 <= io_write_0_data;
      end
      if(_zz_1[27]) begin
        regFile_27 <= io_write_0_data;
      end
      if(_zz_1[28]) begin
        regFile_28 <= io_write_0_data;
      end
      if(_zz_1[29]) begin
        regFile_29 <= io_write_0_data;
      end
      if(_zz_1[30]) begin
        regFile_30 <= io_write_0_data;
      end
      if(_zz_1[31]) begin
        regFile_31 <= io_write_0_data;
      end
      if(_zz_1[32]) begin
        regFile_32 <= io_write_0_data;
      end
      if(_zz_1[33]) begin
        regFile_33 <= io_write_0_data;
      end
      if(_zz_1[34]) begin
        regFile_34 <= io_write_0_data;
      end
      if(_zz_1[35]) begin
        regFile_35 <= io_write_0_data;
      end
      if(_zz_1[36]) begin
        regFile_36 <= io_write_0_data;
      end
      if(_zz_1[37]) begin
        regFile_37 <= io_write_0_data;
      end
      if(_zz_1[38]) begin
        regFile_38 <= io_write_0_data;
      end
      if(_zz_1[39]) begin
        regFile_39 <= io_write_0_data;
      end
      if(_zz_1[40]) begin
        regFile_40 <= io_write_0_data;
      end
      if(_zz_1[41]) begin
        regFile_41 <= io_write_0_data;
      end
      if(_zz_1[42]) begin
        regFile_42 <= io_write_0_data;
      end
      if(_zz_1[43]) begin
        regFile_43 <= io_write_0_data;
      end
      if(_zz_1[44]) begin
        regFile_44 <= io_write_0_data;
      end
      if(_zz_1[45]) begin
        regFile_45 <= io_write_0_data;
      end
      if(_zz_1[46]) begin
        regFile_46 <= io_write_0_data;
      end
      if(_zz_1[47]) begin
        regFile_47 <= io_write_0_data;
      end
      if(_zz_1[48]) begin
        regFile_48 <= io_write_0_data;
      end
      if(_zz_1[49]) begin
        regFile_49 <= io_write_0_data;
      end
      if(_zz_1[50]) begin
        regFile_50 <= io_write_0_data;
      end
      if(_zz_1[51]) begin
        regFile_51 <= io_write_0_data;
      end
      if(_zz_1[52]) begin
        regFile_52 <= io_write_0_data;
      end
      if(_zz_1[53]) begin
        regFile_53 <= io_write_0_data;
      end
      if(_zz_1[54]) begin
        regFile_54 <= io_write_0_data;
      end
      if(_zz_1[55]) begin
        regFile_55 <= io_write_0_data;
      end
      if(_zz_1[56]) begin
        regFile_56 <= io_write_0_data;
      end
      if(_zz_1[57]) begin
        regFile_57 <= io_write_0_data;
      end
      if(_zz_1[58]) begin
        regFile_58 <= io_write_0_data;
      end
      if(_zz_1[59]) begin
        regFile_59 <= io_write_0_data;
      end
      if(_zz_1[60]) begin
        regFile_60 <= io_write_0_data;
      end
      if(_zz_1[61]) begin
        regFile_61 <= io_write_0_data;
      end
      if(_zz_1[62]) begin
        regFile_62 <= io_write_0_data;
      end
      if(_zz_1[63]) begin
        regFile_63 <= io_write_0_data;
      end
    end
    if(when_PRF_l27_1) begin
      if(_zz_2[0]) begin
        regFile_0 <= io_write_1_data;
      end
      if(_zz_2[1]) begin
        regFile_1 <= io_write_1_data;
      end
      if(_zz_2[2]) begin
        regFile_2 <= io_write_1_data;
      end
      if(_zz_2[3]) begin
        regFile_3 <= io_write_1_data;
      end
      if(_zz_2[4]) begin
        regFile_4 <= io_write_1_data;
      end
      if(_zz_2[5]) begin
        regFile_5 <= io_write_1_data;
      end
      if(_zz_2[6]) begin
        regFile_6 <= io_write_1_data;
      end
      if(_zz_2[7]) begin
        regFile_7 <= io_write_1_data;
      end
      if(_zz_2[8]) begin
        regFile_8 <= io_write_1_data;
      end
      if(_zz_2[9]) begin
        regFile_9 <= io_write_1_data;
      end
      if(_zz_2[10]) begin
        regFile_10 <= io_write_1_data;
      end
      if(_zz_2[11]) begin
        regFile_11 <= io_write_1_data;
      end
      if(_zz_2[12]) begin
        regFile_12 <= io_write_1_data;
      end
      if(_zz_2[13]) begin
        regFile_13 <= io_write_1_data;
      end
      if(_zz_2[14]) begin
        regFile_14 <= io_write_1_data;
      end
      if(_zz_2[15]) begin
        regFile_15 <= io_write_1_data;
      end
      if(_zz_2[16]) begin
        regFile_16 <= io_write_1_data;
      end
      if(_zz_2[17]) begin
        regFile_17 <= io_write_1_data;
      end
      if(_zz_2[18]) begin
        regFile_18 <= io_write_1_data;
      end
      if(_zz_2[19]) begin
        regFile_19 <= io_write_1_data;
      end
      if(_zz_2[20]) begin
        regFile_20 <= io_write_1_data;
      end
      if(_zz_2[21]) begin
        regFile_21 <= io_write_1_data;
      end
      if(_zz_2[22]) begin
        regFile_22 <= io_write_1_data;
      end
      if(_zz_2[23]) begin
        regFile_23 <= io_write_1_data;
      end
      if(_zz_2[24]) begin
        regFile_24 <= io_write_1_data;
      end
      if(_zz_2[25]) begin
        regFile_25 <= io_write_1_data;
      end
      if(_zz_2[26]) begin
        regFile_26 <= io_write_1_data;
      end
      if(_zz_2[27]) begin
        regFile_27 <= io_write_1_data;
      end
      if(_zz_2[28]) begin
        regFile_28 <= io_write_1_data;
      end
      if(_zz_2[29]) begin
        regFile_29 <= io_write_1_data;
      end
      if(_zz_2[30]) begin
        regFile_30 <= io_write_1_data;
      end
      if(_zz_2[31]) begin
        regFile_31 <= io_write_1_data;
      end
      if(_zz_2[32]) begin
        regFile_32 <= io_write_1_data;
      end
      if(_zz_2[33]) begin
        regFile_33 <= io_write_1_data;
      end
      if(_zz_2[34]) begin
        regFile_34 <= io_write_1_data;
      end
      if(_zz_2[35]) begin
        regFile_35 <= io_write_1_data;
      end
      if(_zz_2[36]) begin
        regFile_36 <= io_write_1_data;
      end
      if(_zz_2[37]) begin
        regFile_37 <= io_write_1_data;
      end
      if(_zz_2[38]) begin
        regFile_38 <= io_write_1_data;
      end
      if(_zz_2[39]) begin
        regFile_39 <= io_write_1_data;
      end
      if(_zz_2[40]) begin
        regFile_40 <= io_write_1_data;
      end
      if(_zz_2[41]) begin
        regFile_41 <= io_write_1_data;
      end
      if(_zz_2[42]) begin
        regFile_42 <= io_write_1_data;
      end
      if(_zz_2[43]) begin
        regFile_43 <= io_write_1_data;
      end
      if(_zz_2[44]) begin
        regFile_44 <= io_write_1_data;
      end
      if(_zz_2[45]) begin
        regFile_45 <= io_write_1_data;
      end
      if(_zz_2[46]) begin
        regFile_46 <= io_write_1_data;
      end
      if(_zz_2[47]) begin
        regFile_47 <= io_write_1_data;
      end
      if(_zz_2[48]) begin
        regFile_48 <= io_write_1_data;
      end
      if(_zz_2[49]) begin
        regFile_49 <= io_write_1_data;
      end
      if(_zz_2[50]) begin
        regFile_50 <= io_write_1_data;
      end
      if(_zz_2[51]) begin
        regFile_51 <= io_write_1_data;
      end
      if(_zz_2[52]) begin
        regFile_52 <= io_write_1_data;
      end
      if(_zz_2[53]) begin
        regFile_53 <= io_write_1_data;
      end
      if(_zz_2[54]) begin
        regFile_54 <= io_write_1_data;
      end
      if(_zz_2[55]) begin
        regFile_55 <= io_write_1_data;
      end
      if(_zz_2[56]) begin
        regFile_56 <= io_write_1_data;
      end
      if(_zz_2[57]) begin
        regFile_57 <= io_write_1_data;
      end
      if(_zz_2[58]) begin
        regFile_58 <= io_write_1_data;
      end
      if(_zz_2[59]) begin
        regFile_59 <= io_write_1_data;
      end
      if(_zz_2[60]) begin
        regFile_60 <= io_write_1_data;
      end
      if(_zz_2[61]) begin
        regFile_61 <= io_write_1_data;
      end
      if(_zz_2[62]) begin
        regFile_62 <= io_write_1_data;
      end
      if(_zz_2[63]) begin
        regFile_63 <= io_write_1_data;
      end
    end
    if(when_PRF_l27_2) begin
      if(_zz_3[0]) begin
        regFile_0 <= io_write_2_data;
      end
      if(_zz_3[1]) begin
        regFile_1 <= io_write_2_data;
      end
      if(_zz_3[2]) begin
        regFile_2 <= io_write_2_data;
      end
      if(_zz_3[3]) begin
        regFile_3 <= io_write_2_data;
      end
      if(_zz_3[4]) begin
        regFile_4 <= io_write_2_data;
      end
      if(_zz_3[5]) begin
        regFile_5 <= io_write_2_data;
      end
      if(_zz_3[6]) begin
        regFile_6 <= io_write_2_data;
      end
      if(_zz_3[7]) begin
        regFile_7 <= io_write_2_data;
      end
      if(_zz_3[8]) begin
        regFile_8 <= io_write_2_data;
      end
      if(_zz_3[9]) begin
        regFile_9 <= io_write_2_data;
      end
      if(_zz_3[10]) begin
        regFile_10 <= io_write_2_data;
      end
      if(_zz_3[11]) begin
        regFile_11 <= io_write_2_data;
      end
      if(_zz_3[12]) begin
        regFile_12 <= io_write_2_data;
      end
      if(_zz_3[13]) begin
        regFile_13 <= io_write_2_data;
      end
      if(_zz_3[14]) begin
        regFile_14 <= io_write_2_data;
      end
      if(_zz_3[15]) begin
        regFile_15 <= io_write_2_data;
      end
      if(_zz_3[16]) begin
        regFile_16 <= io_write_2_data;
      end
      if(_zz_3[17]) begin
        regFile_17 <= io_write_2_data;
      end
      if(_zz_3[18]) begin
        regFile_18 <= io_write_2_data;
      end
      if(_zz_3[19]) begin
        regFile_19 <= io_write_2_data;
      end
      if(_zz_3[20]) begin
        regFile_20 <= io_write_2_data;
      end
      if(_zz_3[21]) begin
        regFile_21 <= io_write_2_data;
      end
      if(_zz_3[22]) begin
        regFile_22 <= io_write_2_data;
      end
      if(_zz_3[23]) begin
        regFile_23 <= io_write_2_data;
      end
      if(_zz_3[24]) begin
        regFile_24 <= io_write_2_data;
      end
      if(_zz_3[25]) begin
        regFile_25 <= io_write_2_data;
      end
      if(_zz_3[26]) begin
        regFile_26 <= io_write_2_data;
      end
      if(_zz_3[27]) begin
        regFile_27 <= io_write_2_data;
      end
      if(_zz_3[28]) begin
        regFile_28 <= io_write_2_data;
      end
      if(_zz_3[29]) begin
        regFile_29 <= io_write_2_data;
      end
      if(_zz_3[30]) begin
        regFile_30 <= io_write_2_data;
      end
      if(_zz_3[31]) begin
        regFile_31 <= io_write_2_data;
      end
      if(_zz_3[32]) begin
        regFile_32 <= io_write_2_data;
      end
      if(_zz_3[33]) begin
        regFile_33 <= io_write_2_data;
      end
      if(_zz_3[34]) begin
        regFile_34 <= io_write_2_data;
      end
      if(_zz_3[35]) begin
        regFile_35 <= io_write_2_data;
      end
      if(_zz_3[36]) begin
        regFile_36 <= io_write_2_data;
      end
      if(_zz_3[37]) begin
        regFile_37 <= io_write_2_data;
      end
      if(_zz_3[38]) begin
        regFile_38 <= io_write_2_data;
      end
      if(_zz_3[39]) begin
        regFile_39 <= io_write_2_data;
      end
      if(_zz_3[40]) begin
        regFile_40 <= io_write_2_data;
      end
      if(_zz_3[41]) begin
        regFile_41 <= io_write_2_data;
      end
      if(_zz_3[42]) begin
        regFile_42 <= io_write_2_data;
      end
      if(_zz_3[43]) begin
        regFile_43 <= io_write_2_data;
      end
      if(_zz_3[44]) begin
        regFile_44 <= io_write_2_data;
      end
      if(_zz_3[45]) begin
        regFile_45 <= io_write_2_data;
      end
      if(_zz_3[46]) begin
        regFile_46 <= io_write_2_data;
      end
      if(_zz_3[47]) begin
        regFile_47 <= io_write_2_data;
      end
      if(_zz_3[48]) begin
        regFile_48 <= io_write_2_data;
      end
      if(_zz_3[49]) begin
        regFile_49 <= io_write_2_data;
      end
      if(_zz_3[50]) begin
        regFile_50 <= io_write_2_data;
      end
      if(_zz_3[51]) begin
        regFile_51 <= io_write_2_data;
      end
      if(_zz_3[52]) begin
        regFile_52 <= io_write_2_data;
      end
      if(_zz_3[53]) begin
        regFile_53 <= io_write_2_data;
      end
      if(_zz_3[54]) begin
        regFile_54 <= io_write_2_data;
      end
      if(_zz_3[55]) begin
        regFile_55 <= io_write_2_data;
      end
      if(_zz_3[56]) begin
        regFile_56 <= io_write_2_data;
      end
      if(_zz_3[57]) begin
        regFile_57 <= io_write_2_data;
      end
      if(_zz_3[58]) begin
        regFile_58 <= io_write_2_data;
      end
      if(_zz_3[59]) begin
        regFile_59 <= io_write_2_data;
      end
      if(_zz_3[60]) begin
        regFile_60 <= io_write_2_data;
      end
      if(_zz_3[61]) begin
        regFile_61 <= io_write_2_data;
      end
      if(_zz_3[62]) begin
        regFile_62 <= io_write_2_data;
      end
      if(_zz_3[63]) begin
        regFile_63 <= io_write_2_data;
      end
    end
    if(when_PRF_l27_3) begin
      if(_zz_4[0]) begin
        regFile_0 <= io_write_3_data;
      end
      if(_zz_4[1]) begin
        regFile_1 <= io_write_3_data;
      end
      if(_zz_4[2]) begin
        regFile_2 <= io_write_3_data;
      end
      if(_zz_4[3]) begin
        regFile_3 <= io_write_3_data;
      end
      if(_zz_4[4]) begin
        regFile_4 <= io_write_3_data;
      end
      if(_zz_4[5]) begin
        regFile_5 <= io_write_3_data;
      end
      if(_zz_4[6]) begin
        regFile_6 <= io_write_3_data;
      end
      if(_zz_4[7]) begin
        regFile_7 <= io_write_3_data;
      end
      if(_zz_4[8]) begin
        regFile_8 <= io_write_3_data;
      end
      if(_zz_4[9]) begin
        regFile_9 <= io_write_3_data;
      end
      if(_zz_4[10]) begin
        regFile_10 <= io_write_3_data;
      end
      if(_zz_4[11]) begin
        regFile_11 <= io_write_3_data;
      end
      if(_zz_4[12]) begin
        regFile_12 <= io_write_3_data;
      end
      if(_zz_4[13]) begin
        regFile_13 <= io_write_3_data;
      end
      if(_zz_4[14]) begin
        regFile_14 <= io_write_3_data;
      end
      if(_zz_4[15]) begin
        regFile_15 <= io_write_3_data;
      end
      if(_zz_4[16]) begin
        regFile_16 <= io_write_3_data;
      end
      if(_zz_4[17]) begin
        regFile_17 <= io_write_3_data;
      end
      if(_zz_4[18]) begin
        regFile_18 <= io_write_3_data;
      end
      if(_zz_4[19]) begin
        regFile_19 <= io_write_3_data;
      end
      if(_zz_4[20]) begin
        regFile_20 <= io_write_3_data;
      end
      if(_zz_4[21]) begin
        regFile_21 <= io_write_3_data;
      end
      if(_zz_4[22]) begin
        regFile_22 <= io_write_3_data;
      end
      if(_zz_4[23]) begin
        regFile_23 <= io_write_3_data;
      end
      if(_zz_4[24]) begin
        regFile_24 <= io_write_3_data;
      end
      if(_zz_4[25]) begin
        regFile_25 <= io_write_3_data;
      end
      if(_zz_4[26]) begin
        regFile_26 <= io_write_3_data;
      end
      if(_zz_4[27]) begin
        regFile_27 <= io_write_3_data;
      end
      if(_zz_4[28]) begin
        regFile_28 <= io_write_3_data;
      end
      if(_zz_4[29]) begin
        regFile_29 <= io_write_3_data;
      end
      if(_zz_4[30]) begin
        regFile_30 <= io_write_3_data;
      end
      if(_zz_4[31]) begin
        regFile_31 <= io_write_3_data;
      end
      if(_zz_4[32]) begin
        regFile_32 <= io_write_3_data;
      end
      if(_zz_4[33]) begin
        regFile_33 <= io_write_3_data;
      end
      if(_zz_4[34]) begin
        regFile_34 <= io_write_3_data;
      end
      if(_zz_4[35]) begin
        regFile_35 <= io_write_3_data;
      end
      if(_zz_4[36]) begin
        regFile_36 <= io_write_3_data;
      end
      if(_zz_4[37]) begin
        regFile_37 <= io_write_3_data;
      end
      if(_zz_4[38]) begin
        regFile_38 <= io_write_3_data;
      end
      if(_zz_4[39]) begin
        regFile_39 <= io_write_3_data;
      end
      if(_zz_4[40]) begin
        regFile_40 <= io_write_3_data;
      end
      if(_zz_4[41]) begin
        regFile_41 <= io_write_3_data;
      end
      if(_zz_4[42]) begin
        regFile_42 <= io_write_3_data;
      end
      if(_zz_4[43]) begin
        regFile_43 <= io_write_3_data;
      end
      if(_zz_4[44]) begin
        regFile_44 <= io_write_3_data;
      end
      if(_zz_4[45]) begin
        regFile_45 <= io_write_3_data;
      end
      if(_zz_4[46]) begin
        regFile_46 <= io_write_3_data;
      end
      if(_zz_4[47]) begin
        regFile_47 <= io_write_3_data;
      end
      if(_zz_4[48]) begin
        regFile_48 <= io_write_3_data;
      end
      if(_zz_4[49]) begin
        regFile_49 <= io_write_3_data;
      end
      if(_zz_4[50]) begin
        regFile_50 <= io_write_3_data;
      end
      if(_zz_4[51]) begin
        regFile_51 <= io_write_3_data;
      end
      if(_zz_4[52]) begin
        regFile_52 <= io_write_3_data;
      end
      if(_zz_4[53]) begin
        regFile_53 <= io_write_3_data;
      end
      if(_zz_4[54]) begin
        regFile_54 <= io_write_3_data;
      end
      if(_zz_4[55]) begin
        regFile_55 <= io_write_3_data;
      end
      if(_zz_4[56]) begin
        regFile_56 <= io_write_3_data;
      end
      if(_zz_4[57]) begin
        regFile_57 <= io_write_3_data;
      end
      if(_zz_4[58]) begin
        regFile_58 <= io_write_3_data;
      end
      if(_zz_4[59]) begin
        regFile_59 <= io_write_3_data;
      end
      if(_zz_4[60]) begin
        regFile_60 <= io_write_3_data;
      end
      if(_zz_4[61]) begin
        regFile_61 <= io_write_3_data;
      end
      if(_zz_4[62]) begin
        regFile_62 <= io_write_3_data;
      end
      if(_zz_4[63]) begin
        regFile_63 <= io_write_3_data;
      end
    end
    if(when_PRF_l27_4) begin
      if(_zz_5[0]) begin
        regFile_0 <= io_write_4_data;
      end
      if(_zz_5[1]) begin
        regFile_1 <= io_write_4_data;
      end
      if(_zz_5[2]) begin
        regFile_2 <= io_write_4_data;
      end
      if(_zz_5[3]) begin
        regFile_3 <= io_write_4_data;
      end
      if(_zz_5[4]) begin
        regFile_4 <= io_write_4_data;
      end
      if(_zz_5[5]) begin
        regFile_5 <= io_write_4_data;
      end
      if(_zz_5[6]) begin
        regFile_6 <= io_write_4_data;
      end
      if(_zz_5[7]) begin
        regFile_7 <= io_write_4_data;
      end
      if(_zz_5[8]) begin
        regFile_8 <= io_write_4_data;
      end
      if(_zz_5[9]) begin
        regFile_9 <= io_write_4_data;
      end
      if(_zz_5[10]) begin
        regFile_10 <= io_write_4_data;
      end
      if(_zz_5[11]) begin
        regFile_11 <= io_write_4_data;
      end
      if(_zz_5[12]) begin
        regFile_12 <= io_write_4_data;
      end
      if(_zz_5[13]) begin
        regFile_13 <= io_write_4_data;
      end
      if(_zz_5[14]) begin
        regFile_14 <= io_write_4_data;
      end
      if(_zz_5[15]) begin
        regFile_15 <= io_write_4_data;
      end
      if(_zz_5[16]) begin
        regFile_16 <= io_write_4_data;
      end
      if(_zz_5[17]) begin
        regFile_17 <= io_write_4_data;
      end
      if(_zz_5[18]) begin
        regFile_18 <= io_write_4_data;
      end
      if(_zz_5[19]) begin
        regFile_19 <= io_write_4_data;
      end
      if(_zz_5[20]) begin
        regFile_20 <= io_write_4_data;
      end
      if(_zz_5[21]) begin
        regFile_21 <= io_write_4_data;
      end
      if(_zz_5[22]) begin
        regFile_22 <= io_write_4_data;
      end
      if(_zz_5[23]) begin
        regFile_23 <= io_write_4_data;
      end
      if(_zz_5[24]) begin
        regFile_24 <= io_write_4_data;
      end
      if(_zz_5[25]) begin
        regFile_25 <= io_write_4_data;
      end
      if(_zz_5[26]) begin
        regFile_26 <= io_write_4_data;
      end
      if(_zz_5[27]) begin
        regFile_27 <= io_write_4_data;
      end
      if(_zz_5[28]) begin
        regFile_28 <= io_write_4_data;
      end
      if(_zz_5[29]) begin
        regFile_29 <= io_write_4_data;
      end
      if(_zz_5[30]) begin
        regFile_30 <= io_write_4_data;
      end
      if(_zz_5[31]) begin
        regFile_31 <= io_write_4_data;
      end
      if(_zz_5[32]) begin
        regFile_32 <= io_write_4_data;
      end
      if(_zz_5[33]) begin
        regFile_33 <= io_write_4_data;
      end
      if(_zz_5[34]) begin
        regFile_34 <= io_write_4_data;
      end
      if(_zz_5[35]) begin
        regFile_35 <= io_write_4_data;
      end
      if(_zz_5[36]) begin
        regFile_36 <= io_write_4_data;
      end
      if(_zz_5[37]) begin
        regFile_37 <= io_write_4_data;
      end
      if(_zz_5[38]) begin
        regFile_38 <= io_write_4_data;
      end
      if(_zz_5[39]) begin
        regFile_39 <= io_write_4_data;
      end
      if(_zz_5[40]) begin
        regFile_40 <= io_write_4_data;
      end
      if(_zz_5[41]) begin
        regFile_41 <= io_write_4_data;
      end
      if(_zz_5[42]) begin
        regFile_42 <= io_write_4_data;
      end
      if(_zz_5[43]) begin
        regFile_43 <= io_write_4_data;
      end
      if(_zz_5[44]) begin
        regFile_44 <= io_write_4_data;
      end
      if(_zz_5[45]) begin
        regFile_45 <= io_write_4_data;
      end
      if(_zz_5[46]) begin
        regFile_46 <= io_write_4_data;
      end
      if(_zz_5[47]) begin
        regFile_47 <= io_write_4_data;
      end
      if(_zz_5[48]) begin
        regFile_48 <= io_write_4_data;
      end
      if(_zz_5[49]) begin
        regFile_49 <= io_write_4_data;
      end
      if(_zz_5[50]) begin
        regFile_50 <= io_write_4_data;
      end
      if(_zz_5[51]) begin
        regFile_51 <= io_write_4_data;
      end
      if(_zz_5[52]) begin
        regFile_52 <= io_write_4_data;
      end
      if(_zz_5[53]) begin
        regFile_53 <= io_write_4_data;
      end
      if(_zz_5[54]) begin
        regFile_54 <= io_write_4_data;
      end
      if(_zz_5[55]) begin
        regFile_55 <= io_write_4_data;
      end
      if(_zz_5[56]) begin
        regFile_56 <= io_write_4_data;
      end
      if(_zz_5[57]) begin
        regFile_57 <= io_write_4_data;
      end
      if(_zz_5[58]) begin
        regFile_58 <= io_write_4_data;
      end
      if(_zz_5[59]) begin
        regFile_59 <= io_write_4_data;
      end
      if(_zz_5[60]) begin
        regFile_60 <= io_write_4_data;
      end
      if(_zz_5[61]) begin
        regFile_61 <= io_write_4_data;
      end
      if(_zz_5[62]) begin
        regFile_62 <= io_write_4_data;
      end
      if(_zz_5[63]) begin
        regFile_63 <= io_write_4_data;
      end
    end
    io_debugRegs_0 <= regFile_0;
    io_debugRegs_1 <= regFile_1;
    io_debugRegs_2 <= regFile_2;
    io_debugRegs_3 <= regFile_3;
    io_debugRegs_4 <= regFile_4;
    io_debugRegs_5 <= regFile_5;
    io_debugRegs_6 <= regFile_6;
    io_debugRegs_7 <= regFile_7;
    io_debugRegs_8 <= regFile_8;
    io_debugRegs_9 <= regFile_9;
    io_debugRegs_10 <= regFile_10;
    io_debugRegs_11 <= regFile_11;
    io_debugRegs_12 <= regFile_12;
    io_debugRegs_13 <= regFile_13;
    io_debugRegs_14 <= regFile_14;
    io_debugRegs_15 <= regFile_15;
    io_debugRegs_16 <= regFile_16;
    io_debugRegs_17 <= regFile_17;
    io_debugRegs_18 <= regFile_18;
    io_debugRegs_19 <= regFile_19;
    io_debugRegs_20 <= regFile_20;
    io_debugRegs_21 <= regFile_21;
    io_debugRegs_22 <= regFile_22;
    io_debugRegs_23 <= regFile_23;
    io_debugRegs_24 <= regFile_24;
    io_debugRegs_25 <= regFile_25;
    io_debugRegs_26 <= regFile_26;
    io_debugRegs_27 <= regFile_27;
    io_debugRegs_28 <= regFile_28;
    io_debugRegs_29 <= regFile_29;
    io_debugRegs_30 <= regFile_30;
    io_debugRegs_31 <= regFile_31;
    io_debugRegs_32 <= regFile_32;
    io_debugRegs_33 <= regFile_33;
    io_debugRegs_34 <= regFile_34;
    io_debugRegs_35 <= regFile_35;
    io_debugRegs_36 <= regFile_36;
    io_debugRegs_37 <= regFile_37;
    io_debugRegs_38 <= regFile_38;
    io_debugRegs_39 <= regFile_39;
    io_debugRegs_40 <= regFile_40;
    io_debugRegs_41 <= regFile_41;
    io_debugRegs_42 <= regFile_42;
    io_debugRegs_43 <= regFile_43;
    io_debugRegs_44 <= regFile_44;
    io_debugRegs_45 <= regFile_45;
    io_debugRegs_46 <= regFile_46;
    io_debugRegs_47 <= regFile_47;
    io_debugRegs_48 <= regFile_48;
    io_debugRegs_49 <= regFile_49;
    io_debugRegs_50 <= regFile_50;
    io_debugRegs_51 <= regFile_51;
    io_debugRegs_52 <= regFile_52;
    io_debugRegs_53 <= regFile_53;
    io_debugRegs_54 <= regFile_54;
    io_debugRegs_55 <= regFile_55;
    io_debugRegs_56 <= regFile_56;
    io_debugRegs_57 <= regFile_57;
    io_debugRegs_58 <= regFile_58;
    io_debugRegs_59 <= regFile_59;
    io_debugRegs_60 <= regFile_60;
    io_debugRegs_61 <= regFile_61;
    io_debugRegs_62 <= regFile_62;
    io_debugRegs_63 <= regFile_63;
  end


endmodule

module DCache (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [31:0]   io_input_payload_src1,
  input  wire [31:0]   io_input_payload_src2,
  input  wire [31:0]   io_input_payload_src3,
  input  wire [4:0]    io_input_payload_robIdx,
  input  wire [31:0]   io_input_payload_branchResult_targetPC,
  input  wire          io_input_payload_branchResult_branchResult,
  input  wire          io_input_payload_branchResult_predictFail,
  input  wire          io_input_payload_exceptionInfo_exception,
  input  wire [5:0]    io_input_payload_exceptionInfo_eCode,
  input  wire [0:0]    io_input_payload_exceptionInfo_eSubCode,
  input  wire [31:0]   io_input_payload_pc,
  input  wire [5:0]    io_input_payload_prd,
  input  wire [3:0]    io_input_payload_uop_lsuOp,
  input  wire [4:0]    io_input_payload_uop_lsuCoOp,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [4:0]    io_output_payload_robIdx,
  output wire [31:0]   io_output_payload_data,
  output wire [5:0]    io_output_payload_prd,
  output wire [31:0]   io_output_payload_branchResult_targetPC,
  output wire          io_output_payload_branchResult_branchResult,
  output wire          io_output_payload_branchResult_predictFail,
  output wire          io_output_payload_exceptionInfo_exception,
  output wire [5:0]    io_output_payload_exceptionInfo_eCode,
  output wire [0:0]    io_output_payload_exceptionInfo_eSubCode,
  output wire          io_wakeOut_0_valid,
  output wire [5:0]    io_wakeOut_0_payload,
  output wire          io_wakeOut_1_valid,
  output wire [5:0]    io_wakeOut_1_payload,
  input  wire [4:0]    io_retireComm_robIdx_0,
  input  wire [4:0]    io_retireComm_robIdx_1,
  input  wire          io_retireComm_allowRetire_0,
  input  wire          io_retireComm_allowRetire_1,
  input  wire          io_tlb_hit,
  input  wire [19:0]   io_tlb_pageInfo_ppn,
  input  wire [1:0]    io_tlb_pageInfo_plv,
  input  wire [1:0]    io_tlb_pageInfo_mat,
  input  wire          io_tlb_pageInfo_d,
  input  wire          io_tlb_pageInfo_v,
  output wire [19:0]   io_tlb_virtPageNumber,
  input  wire [1:0]    _zz_when_LSU_l217,
  input  wire [31:0]   io_llBitComm_actualAddr,
  output wire [31:0]   io_llBitComm_toUpdateAddr,
  output wire          io_llBitComm_wen,
  input  wire          _zz_scMatchHit,
  output wire          io_ctrl_busy,
  input  wire          io_ctrl_stall,
  input  wire [31:0]   io_ctrl_cacopVA,
  input  wire          io_ctrl_cacopStoreTag,
  input  wire          io_ctrl_cacopIndexInvalidate,
  input  wire          io_ctrl_cacopHitInvalidate,
  output wire          io_specialOpBufferUpdate_valid,
  output wire [3:0]    io_specialOpBufferUpdate_payload_uop_lsuOp,
  output wire [4:0]    io_specialOpBufferUpdate_payload_uop_lsuCoOp,
  output wire [31:0]   io_specialOpBufferUpdate_payload_vaddr,
  output wire [9:0]    io_specialOpBufferUpdate_payload_asid,
  input  wire          io_flush,
  output wire [4:0]    io_badv_robIdx,
  output wire [31:0]   io_badv_vaddr,
  output wire          io_badv_wen,
  output wire [3:0]    io_axi_arid,
  output wire [31:0]   io_axi_araddr,
  output wire [7:0]    io_axi_arlen,
  output wire [2:0]    io_axi_arsize,
  output wire [1:0]    io_axi_arburst,
  output wire [1:0]    io_axi_arlock,
  output wire [3:0]    io_axi_arcache,
  output wire [2:0]    io_axi_arprot,
  output reg           io_axi_arvalid,
  input  wire          io_axi_arready,
  input  wire [3:0]    io_axi_rid,
  input  wire [31:0]   io_axi_rdata,
  input  wire [1:0]    io_axi_rresp,
  input  wire          io_axi_rlast,
  input  wire          io_axi_rvalid,
  output reg           io_axi_rready,
  output wire [3:0]    io_axi_awid,
  output wire [31:0]   io_axi_awaddr,
  output wire [7:0]    io_axi_awlen,
  output wire [2:0]    io_axi_awsize,
  output wire [1:0]    io_axi_awburst,
  output wire [1:0]    io_axi_awlock,
  output wire [3:0]    io_axi_awcache,
  output wire [2:0]    io_axi_awprot,
  output reg           io_axi_awvalid,
  input  wire          io_axi_awready,
  output wire [3:0]    io_axi_wid,
  output wire [31:0]   io_axi_wdata,
  output wire [3:0]    io_axi_wstrb,
  output wire          io_axi_wlast,
  output reg           io_axi_wvalid,
  input  wire          io_axi_wready,
  input  wire [3:0]    io_axi_bid,
  input  wire [1:0]    io_axi_bresp,
  input  wire          io_axi_bvalid,
  output wire          io_axi_bready,
  output wire [31:0]   io_storeData,
  output wire [3:0]    io_storeMask,
  output wire [3:0]    io_loadMask,
  output wire [31:0]   io_VAddr,
  output wire [31:0]   io_PAddr,
  input  wire          aclk,
  input  wire          aresetn
);
  localparam LSUOp_cacop = 4'd0;
  localparam LSUOp_tlbsrch = 4'd1;
  localparam LSUOp_tlbrd = 4'd2;
  localparam LSUOp_tlbwr = 4'd3;
  localparam LSUOp_tlbfill = 4'd4;
  localparam LSUOp_invtlb = 4'd5;
  localparam LSUOp_ll = 4'd6;
  localparam LSUOp_sc = 4'd7;
  localparam LSUOp_ld = 4'd8;
  localparam LSUOp_ldu = 4'd9;
  localparam LSUOp_st = 4'd10;
  localparam LSUOp_preld = 4'd11;
  localparam LSUOp_dbar = 4'd12;
  localparam LSUOp_ibar = 4'd13;
  localparam LSUSizeOp_byte_1 = 4'd1;
  localparam LSUSizeOp_halfword = 4'd3;
  localparam LSUSizeOp_word = 4'd15;
  localparam axiCtrl_enumDef_BOOT = 3'd0;
  localparam axiCtrl_enumDef_idle = 3'd1;
  localparam axiCtrl_enumDef_readReq = 3'd2;
  localparam axiCtrl_enumDef_readFirst = 3'd3;
  localparam axiCtrl_enumDef_read = 3'd4;
  localparam axiCtrl_enumDef_writeReq = 3'd5;
  localparam axiCtrl_enumDef_write = 3'd6;
  localparam rollbackCtrl_enumDef_BOOT = 2'd0;
  localparam rollbackCtrl_enumDef_idle = 2'd1;
  localparam rollbackCtrl_enumDef_rollback = 2'd2;

  wire                data_0_portA_en;
  wire                data_0_portB_en;
  wire                data_1_portA_en;
  wire                data_1_portB_en;
  wire                data_2_portA_en;
  wire                data_2_portB_en;
  wire                data_3_portA_en;
  wire                data_3_portB_en;
  wire                tag_0_wr_en;
  wire       [0:0]    tag_0_wr_mask;
  wire       [4:0]    tag_0_wr_addr;
  wire       [20:0]   tag_0_wr_data;
  wire                tag_0_rd_en;
  wire       [4:0]    tag_0_rd_addr;
  wire                tag_1_wr_en;
  wire       [0:0]    tag_1_wr_mask;
  wire       [4:0]    tag_1_wr_addr;
  wire       [20:0]   tag_1_wr_data;
  wire                tag_1_rd_en;
  wire       [4:0]    tag_1_rd_addr;
  wire                tag_2_wr_en;
  wire       [0:0]    tag_2_wr_mask;
  wire       [4:0]    tag_2_wr_addr;
  wire       [20:0]   tag_2_wr_data;
  wire                tag_2_rd_en;
  wire       [4:0]    tag_2_rd_addr;
  wire                tag_3_wr_en;
  wire       [0:0]    tag_3_wr_mask;
  wire       [4:0]    tag_3_wr_addr;
  wire       [20:0]   tag_3_wr_data;
  wire                tag_3_rd_en;
  wire       [4:0]    tag_3_rd_addr;
  wire       [31:0]   data_0_portA_rdData;
  wire       [31:0]   data_0_portB_rdData;
  wire       [31:0]   data_1_portA_rdData;
  wire       [31:0]   data_1_portB_rdData;
  wire       [31:0]   data_2_portA_rdData;
  wire       [31:0]   data_2_portB_rdData;
  wire       [31:0]   data_3_portA_rdData;
  wire       [31:0]   data_3_portB_rdData;
  wire       [20:0]   tag_0_rd_data;
  wire       [20:0]   tag_1_rd_data;
  wire       [20:0]   tag_2_rd_data;
  wire       [20:0]   tag_3_rd_data;
  wire       [31:0]   _zz_stage1Out_payload_storeData;
  wire       [0:0]    _zz_stage1Out_payload_lsCtrlBundle_size;
  wire       [1:0]    _zz_stage1Out_payload_lsCtrlBundle_size_1;
  wire       [1:0]    _zz_stage1Out_payload_lsCtrlBundle_size_2;
  wire       [4:0]    _zz_stage1Out_payload_checkTLBException;
  wire       [1:0]    _zz_stage1Out_payload_checkTLBException_1;
  wire       [31:0]   _zz_portAddr0;
  wire       [31:0]   _zz_portAddr1;
  wire       [31:0]   _zz_portAddr1_1;
  reg                 _zz_stage1Out_payload_wayValid;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_1;
  wire       [31:0]   _zz_stage1Out_payload_wayValid_2;
  reg                 _zz_stage1Out_payload_wayDirty;
  wire       [4:0]    _zz_stage1Out_payload_wayDirty_1;
  wire       [31:0]   _zz_stage1Out_payload_wayDirty_2;
  wire       [1:0]    _zz_hit;
  wire       [0:0]    _zz_hit_1;
  reg                 _zz_stage1Out_payload_wayValid_3;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_4;
  wire       [31:0]   _zz_stage1Out_payload_wayValid_5;
  reg                 _zz_stage1Out_payload_wayDirty_3;
  wire       [4:0]    _zz_stage1Out_payload_wayDirty_4;
  wire       [31:0]   _zz_stage1Out_payload_wayDirty_5;
  wire       [1:0]    _zz_hit_2;
  wire       [0:0]    _zz_hit_3;
  reg                 _zz_stage1Out_payload_wayValid_6;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_7;
  wire       [31:0]   _zz_stage1Out_payload_wayValid_8;
  reg                 _zz_stage1Out_payload_wayDirty_6;
  wire       [4:0]    _zz_stage1Out_payload_wayDirty_7;
  wire       [31:0]   _zz_stage1Out_payload_wayDirty_8;
  wire       [1:0]    _zz_hit_4;
  wire       [0:0]    _zz_hit_5;
  reg                 _zz_stage1Out_payload_wayValid_9;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_10;
  wire       [31:0]   _zz_stage1Out_payload_wayValid_11;
  reg                 _zz_stage1Out_payload_wayDirty_9;
  wire       [4:0]    _zz_stage1Out_payload_wayDirty_10;
  wire       [31:0]   _zz_stage1Out_payload_wayDirty_11;
  wire       [1:0]    _zz_hit_6;
  wire       [0:0]    _zz_hit_7;
  wire       [3:0]    _zz_exceptionInfo1_eCode;
  wire       [3:0]    _zz_exceptionInfo1_eCode_1;
  wire       [5:0]    _zz_exceptionInfo2_eCode;
  wire       [0:0]    _zz_exceptionInfo2_eCode_1;
  wire       [5:0]    _zz_exceptionInfo2_eCode_2;
  wire       [1:0]    _zz_exceptionInfo2_eCode_3;
  wire       [2:0]    _zz_exceptionInfo2_eCode_4;
  wire       [2:0]    _zz_exceptionInfo2_eCode_5;
  wire       [2:0]    _zz_exceptionInfo2_eCode_6;
  wire       [2:0]    _zz_writeBufferHeadNext_8;
  wire       [3:0]    _zz_writeBufferHeadNext_9;
  wire       [3:0]    _zz_writeBufferHeadNext_10;
  reg        [3:0]    _zz_writeBufferHeadNext_11;
  wire       [2:0]    _zz_writeBufferHeadNext_12;
  reg        [3:0]    _zz_writeBufferHeadNext_13;
  wire       [2:0]    _zz_writeBufferHeadNext_14;
  reg        [3:0]    _zz_writeBufferHeadNext_15;
  wire       [2:0]    _zz_writeBufferHeadNext_16;
  wire       [1:0]    _zz_writeBufferHeadNext_17;
  reg                 _zz__zz_writeBufferAvail;
  reg        [4:0]    _zz_latestWrite_robIdx;
  reg        [3:0]    _zz_latestWrite_waySelect;
  reg        [31:0]   _zz_latestWrite_prevData;
  reg                 _zz_latestWrite_prevDirty;
  reg        [8:0]    _zz_latestWrite_index;
  reg                 _zz_latestWrite_miss;
  wire       [1:0]    _zz_writeBufferAppend;
  wire       [0:0]    _zz_writeBufferAppend_1;
  reg        [31:0]   _zz__zz_writeBuffer_0_prevData;
  reg                 _zz__zz_writeBuffer_0_prevDirty;
  wire       [0:0]    _zz__zz_19;
  reg                 _zz_missBuffer_0_writeBack_8;
  reg        [20:0]   _zz_missBuffer_0_prevPaddr;
  wire       [1:0]    _zz_when_LSU_l335;
  wire       [0:0]    _zz_when_LSU_l335_1;
  wire       [1:0]    _zz_dirtyUpdate;
  wire       [0:0]    _zz_dirtyUpdate_1;
  wire       [31:0]   _zz__zz_53;
  wire       [31:0]   _zz__zz_54;
  wire       [31:0]   _zz__zz_55;
  wire       [31:0]   _zz__zz_56;
  wire       [31:0]   _zz_when_LSU_l357;
  wire       [31:0]   _zz_when_LSU_l357_1;
  wire       [0:0]    _zz_io_axi_arid;
  wire       [7:0]    _zz_io_axi_arlen;
  wire       [3:0]    _zz_io_axi_arlen_1;
  wire       [2:0]    _zz_io_axi_arsize;
  wire       [1:0]    _zz_io_axi_arsize_1;
  wire       [0:0]    _zz_io_axi_awid;
  wire       [3:0]    _zz_io_axi_awlen;
  wire       [2:0]    _zz_io_axi_awsize;
  wire       [1:0]    _zz_io_axi_awsize_1;
  wire       [0:0]    _zz_io_axi_awburst;
  wire       [0:0]    _zz_io_axi_wid;
  reg        [31:0]   _zz_io_axi_wdata_2;
  wire       [1:0]    _zz_io_axi_wdata_3;
  wire       [1:0]    _zz__zz_missBufferAllowMask;
  wire       [8:0]    _zz__zz_missBufferPreAllowMask;
  wire       [4:0]    _zz__zz_missBufferPreAllowMask_1;
  wire       [8:0]    _zz__zz_missBufferPreAllowMask_2;
  wire       [4:0]    _zz__zz_missBufferPreAllowMask_3;
  wire       [8:0]    _zz__zz_missBufferPreAllowMask_4;
  wire       [4:0]    _zz__zz_missBufferPreAllowMask_5;
  wire       [8:0]    _zz__zz_missBufferPreAllowMask_6;
  wire       [4:0]    _zz__zz_missBufferPreAllowMask_7;
  wire       [8:0]    _zz__zz_missBufferPreAllowMask_8;
  wire       [4:0]    _zz__zz_missBufferPreAllowMask_9;
  wire       [8:0]    _zz__zz_missBufferPreAllowMask_10;
  wire       [4:0]    _zz__zz_missBufferPreAllowMask_11;
  wire       [8:0]    _zz__zz_missBufferPreAllowMask_12;
  wire       [4:0]    _zz__zz_missBufferPreAllowMask_13;
  wire       [8:0]    _zz__zz_missBufferPreAllowMask_14;
  wire       [4:0]    _zz__zz_missBufferPreAllowMask_15;
  reg        [20:0]   _zz_cacopPAddr;
  wire       [1:0]    _zz_cacopPAddr_1;
  reg                 _zz__zz_wayToReplace;
  wire       [4:0]    _zz__zz_wayToReplace_1;
  reg                 _zz__zz_wayToReplace_2;
  wire       [4:0]    _zz__zz_wayToReplace_3;
  reg                 _zz__zz_wayToReplace_1_1;
  wire       [4:0]    _zz__zz_wayToReplace_1_2;
  reg                 _zz__zz_wayToReplace_1_3;
  wire       [4:0]    _zz__zz_wayToReplace_1_4;
  reg                 _zz__zz_wayToReplace_2_1;
  wire       [4:0]    _zz__zz_wayToReplace_2_2;
  reg                 _zz__zz_wayToReplace_2_3;
  wire       [4:0]    _zz__zz_wayToReplace_2_4;
  reg                 _zz__zz_wayToReplace_3_1;
  wire       [4:0]    _zz__zz_wayToReplace_3_2;
  reg                 _zz__zz_wayToReplace_3_3;
  wire       [4:0]    _zz__zz_wayToReplace_3_4;
  wire       [0:0]    _zz_dataShuffle_0_3;
  wire       [13:0]   _zz_dataShuffle_0_4;
  wire       [0:0]    _zz_dataShuffle_0_5;
  wire       [5:0]    _zz_dataShuffle_0_6;
  wire       [0:0]    _zz_dataShuffle_1_3;
  wire       [13:0]   _zz_dataShuffle_1_4;
  wire       [0:0]    _zz_dataShuffle_1_5;
  wire       [5:0]    _zz_dataShuffle_1_6;
  wire       [0:0]    _zz_dataShuffle_2_3;
  wire       [13:0]   _zz_dataShuffle_2_4;
  wire       [0:0]    _zz_dataShuffle_2_5;
  wire       [5:0]    _zz_dataShuffle_2_6;
  wire       [0:0]    _zz_dataShuffle_3_3;
  wire       [13:0]   _zz_dataShuffle_3_4;
  wire       [0:0]    _zz_dataShuffle_3_5;
  wire       [5:0]    _zz_dataShuffle_3_6;
  wire       [0:0]    _zz_axiShuffle_2;
  wire       [13:0]   _zz_axiShuffle_3;
  wire       [0:0]    _zz_axiShuffle_4;
  wire       [5:0]    _zz_axiShuffle_5;
  reg        [31:0]   _zz_io_output_payload_data_3;
  wire       [3:0]    _zz_cacopWay;
  wire       [31:0]   _zz__zz_65;
  wire       [31:0]   _zz__zz_66;
  wire       [31:0]   _zz__zz_67;
  wire       [31:0]   _zz__zz_68;
  wire       [31:0]   _zz__zz_69;
  wire       [31:0]   _zz__zz_70;
  wire       [31:0]   _zz__zz_71;
  wire       [31:0]   _zz__zz_72;
  wire       [3:0]    _zz_transferRAddrMid;
  wire       [3:0]    _zz_transferRAddrMid_1;
  wire       [3:0]    _zz_transferWAddrMid;
  reg                 _zz_when_LSU_l567;
  wire       [31:0]   _zz_wr_addr;
  wire       [31:0]   _zz_wr_data;
  wire       [31:0]   _zz_rd_addr;
  wire       [31:0]   _zz_wr_addr_1;
  wire       [31:0]   _zz_wr_data_1;
  wire       [31:0]   _zz_rd_addr_1;
  wire       [31:0]   _zz_wr_addr_2;
  wire       [31:0]   _zz_wr_data_2;
  wire       [31:0]   _zz_rd_addr_2;
  wire       [31:0]   _zz_wr_addr_3;
  wire       [31:0]   _zz_wr_data_3;
  wire       [31:0]   _zz_rd_addr_3;
  reg                 _zz_wr_en;
  reg                 _zz_wr_en_1;
  reg                 _zz_wr_en_2;
  reg                 _zz_wr_en_3;
  wire       [31:0]   address;
  reg                 valid_0_0;
  reg                 valid_0_1;
  reg                 valid_0_2;
  reg                 valid_0_3;
  reg                 valid_0_4;
  reg                 valid_0_5;
  reg                 valid_0_6;
  reg                 valid_0_7;
  reg                 valid_0_8;
  reg                 valid_0_9;
  reg                 valid_0_10;
  reg                 valid_0_11;
  reg                 valid_0_12;
  reg                 valid_0_13;
  reg                 valid_0_14;
  reg                 valid_0_15;
  reg                 valid_0_16;
  reg                 valid_0_17;
  reg                 valid_0_18;
  reg                 valid_0_19;
  reg                 valid_0_20;
  reg                 valid_0_21;
  reg                 valid_0_22;
  reg                 valid_0_23;
  reg                 valid_0_24;
  reg                 valid_0_25;
  reg                 valid_0_26;
  reg                 valid_0_27;
  reg                 valid_0_28;
  reg                 valid_0_29;
  reg                 valid_0_30;
  reg                 valid_0_31;
  reg                 valid_1_0;
  reg                 valid_1_1;
  reg                 valid_1_2;
  reg                 valid_1_3;
  reg                 valid_1_4;
  reg                 valid_1_5;
  reg                 valid_1_6;
  reg                 valid_1_7;
  reg                 valid_1_8;
  reg                 valid_1_9;
  reg                 valid_1_10;
  reg                 valid_1_11;
  reg                 valid_1_12;
  reg                 valid_1_13;
  reg                 valid_1_14;
  reg                 valid_1_15;
  reg                 valid_1_16;
  reg                 valid_1_17;
  reg                 valid_1_18;
  reg                 valid_1_19;
  reg                 valid_1_20;
  reg                 valid_1_21;
  reg                 valid_1_22;
  reg                 valid_1_23;
  reg                 valid_1_24;
  reg                 valid_1_25;
  reg                 valid_1_26;
  reg                 valid_1_27;
  reg                 valid_1_28;
  reg                 valid_1_29;
  reg                 valid_1_30;
  reg                 valid_1_31;
  reg                 valid_2_0;
  reg                 valid_2_1;
  reg                 valid_2_2;
  reg                 valid_2_3;
  reg                 valid_2_4;
  reg                 valid_2_5;
  reg                 valid_2_6;
  reg                 valid_2_7;
  reg                 valid_2_8;
  reg                 valid_2_9;
  reg                 valid_2_10;
  reg                 valid_2_11;
  reg                 valid_2_12;
  reg                 valid_2_13;
  reg                 valid_2_14;
  reg                 valid_2_15;
  reg                 valid_2_16;
  reg                 valid_2_17;
  reg                 valid_2_18;
  reg                 valid_2_19;
  reg                 valid_2_20;
  reg                 valid_2_21;
  reg                 valid_2_22;
  reg                 valid_2_23;
  reg                 valid_2_24;
  reg                 valid_2_25;
  reg                 valid_2_26;
  reg                 valid_2_27;
  reg                 valid_2_28;
  reg                 valid_2_29;
  reg                 valid_2_30;
  reg                 valid_2_31;
  reg                 valid_3_0;
  reg                 valid_3_1;
  reg                 valid_3_2;
  reg                 valid_3_3;
  reg                 valid_3_4;
  reg                 valid_3_5;
  reg                 valid_3_6;
  reg                 valid_3_7;
  reg                 valid_3_8;
  reg                 valid_3_9;
  reg                 valid_3_10;
  reg                 valid_3_11;
  reg                 valid_3_12;
  reg                 valid_3_13;
  reg                 valid_3_14;
  reg                 valid_3_15;
  reg                 valid_3_16;
  reg                 valid_3_17;
  reg                 valid_3_18;
  reg                 valid_3_19;
  reg                 valid_3_20;
  reg                 valid_3_21;
  reg                 valid_3_22;
  reg                 valid_3_23;
  reg                 valid_3_24;
  reg                 valid_3_25;
  reg                 valid_3_26;
  reg                 valid_3_27;
  reg                 valid_3_28;
  reg                 valid_3_29;
  reg                 valid_3_30;
  reg                 valid_3_31;
  reg                 dirty_0_0;
  reg                 dirty_0_1;
  reg                 dirty_0_2;
  reg                 dirty_0_3;
  reg                 dirty_0_4;
  reg                 dirty_0_5;
  reg                 dirty_0_6;
  reg                 dirty_0_7;
  reg                 dirty_0_8;
  reg                 dirty_0_9;
  reg                 dirty_0_10;
  reg                 dirty_0_11;
  reg                 dirty_0_12;
  reg                 dirty_0_13;
  reg                 dirty_0_14;
  reg                 dirty_0_15;
  reg                 dirty_0_16;
  reg                 dirty_0_17;
  reg                 dirty_0_18;
  reg                 dirty_0_19;
  reg                 dirty_0_20;
  reg                 dirty_0_21;
  reg                 dirty_0_22;
  reg                 dirty_0_23;
  reg                 dirty_0_24;
  reg                 dirty_0_25;
  reg                 dirty_0_26;
  reg                 dirty_0_27;
  reg                 dirty_0_28;
  reg                 dirty_0_29;
  reg                 dirty_0_30;
  reg                 dirty_0_31;
  reg                 dirty_1_0;
  reg                 dirty_1_1;
  reg                 dirty_1_2;
  reg                 dirty_1_3;
  reg                 dirty_1_4;
  reg                 dirty_1_5;
  reg                 dirty_1_6;
  reg                 dirty_1_7;
  reg                 dirty_1_8;
  reg                 dirty_1_9;
  reg                 dirty_1_10;
  reg                 dirty_1_11;
  reg                 dirty_1_12;
  reg                 dirty_1_13;
  reg                 dirty_1_14;
  reg                 dirty_1_15;
  reg                 dirty_1_16;
  reg                 dirty_1_17;
  reg                 dirty_1_18;
  reg                 dirty_1_19;
  reg                 dirty_1_20;
  reg                 dirty_1_21;
  reg                 dirty_1_22;
  reg                 dirty_1_23;
  reg                 dirty_1_24;
  reg                 dirty_1_25;
  reg                 dirty_1_26;
  reg                 dirty_1_27;
  reg                 dirty_1_28;
  reg                 dirty_1_29;
  reg                 dirty_1_30;
  reg                 dirty_1_31;
  reg                 dirty_2_0;
  reg                 dirty_2_1;
  reg                 dirty_2_2;
  reg                 dirty_2_3;
  reg                 dirty_2_4;
  reg                 dirty_2_5;
  reg                 dirty_2_6;
  reg                 dirty_2_7;
  reg                 dirty_2_8;
  reg                 dirty_2_9;
  reg                 dirty_2_10;
  reg                 dirty_2_11;
  reg                 dirty_2_12;
  reg                 dirty_2_13;
  reg                 dirty_2_14;
  reg                 dirty_2_15;
  reg                 dirty_2_16;
  reg                 dirty_2_17;
  reg                 dirty_2_18;
  reg                 dirty_2_19;
  reg                 dirty_2_20;
  reg                 dirty_2_21;
  reg                 dirty_2_22;
  reg                 dirty_2_23;
  reg                 dirty_2_24;
  reg                 dirty_2_25;
  reg                 dirty_2_26;
  reg                 dirty_2_27;
  reg                 dirty_2_28;
  reg                 dirty_2_29;
  reg                 dirty_2_30;
  reg                 dirty_2_31;
  reg                 dirty_3_0;
  reg                 dirty_3_1;
  reg                 dirty_3_2;
  reg                 dirty_3_3;
  reg                 dirty_3_4;
  reg                 dirty_3_5;
  reg                 dirty_3_6;
  reg                 dirty_3_7;
  reg                 dirty_3_8;
  reg                 dirty_3_9;
  reg                 dirty_3_10;
  reg                 dirty_3_11;
  reg                 dirty_3_12;
  reg                 dirty_3_13;
  reg                 dirty_3_14;
  reg                 dirty_3_15;
  reg                 dirty_3_16;
  reg                 dirty_3_17;
  reg                 dirty_3_18;
  reg                 dirty_3_19;
  reg                 dirty_3_20;
  reg                 dirty_3_21;
  reg                 dirty_3_22;
  reg                 dirty_3_23;
  reg                 dirty_3_24;
  reg                 dirty_3_25;
  reg                 dirty_3_26;
  reg                 dirty_3_27;
  reg                 dirty_3_28;
  reg                 dirty_3_29;
  reg                 dirty_3_30;
  reg                 dirty_3_31;
  wire       [31:0]   dataRead_0;
  wire       [31:0]   dataRead_1;
  wire       [31:0]   dataRead_2;
  wire       [31:0]   dataRead_3;
  wire       [20:0]   tagRead_0;
  wire       [20:0]   tagRead_1;
  wire       [20:0]   tagRead_2;
  wire       [20:0]   tagRead_3;
  reg        [3:0]    hit;
  wire                miss;
  wire                missBufferAvail;
  reg        [3:0]    wayToReplace;
  wire       [3:0]    realLSMask;
  wire                stall;
  wire                cacopActive;
  wire                cacopEn;
  reg                 rollingBack;
  wire                writeBufferAvail;
  wire                writeBufferAppend;
  reg                 writeBufferUpdate;
  reg                 refilling;
  wire                exceptionInfo_exception;
  wire       [5:0]    exceptionInfo_eCode;
  wire       [0:0]    exceptionInfo_eSubCode;
  reg                 exceptionInfo1_exception;
  reg        [5:0]    exceptionInfo1_eCode;
  reg        [0:0]    exceptionInfo1_eSubCode;
  reg                 exceptionInfo2_exception;
  reg        [5:0]    exceptionInfo2_eCode;
  reg        [0:0]    exceptionInfo2_eSubCode;
  wire       [3:0]    wayDirty;
  reg        [3:0]    wayDirtyBypass;
  wire                stage1Out_valid;
  reg                 stage1Out_ready;
  wire       [4:0]    stage1Out_payload_robIdx;
  wire       [5:0]    stage1Out_payload_prd;
  wire       [31:0]   stage1Out_payload_branchResult_targetPC;
  wire                stage1Out_payload_branchResult_branchResult;
  wire                stage1Out_payload_branchResult_predictFail;
  wire                stage1Out_payload_exceptionInfo_exception;
  wire       [5:0]    stage1Out_payload_exceptionInfo_eCode;
  wire       [0:0]    stage1Out_payload_exceptionInfo_eSubCode;
  wire       [31:0]   stage1Out_payload_storeData;
  wire                stage1Out_payload_lsCtrlBundle_load;
  wire                stage1Out_payload_lsCtrlBundle_store;
  wire                stage1Out_payload_lsCtrlBundle_signed;
  wire                stage1Out_payload_lsCtrlBundle_ll;
  wire                stage1Out_payload_lsCtrlBundle_sc;
  wire       [3:0]    stage1Out_payload_lsCtrlBundle_lsMask;
  reg        [2:0]    stage1Out_payload_lsCtrlBundle_size;
  wire                stage1Out_payload_lsCtrlBundle_normalMemOp;
  wire       [31:0]   stage1Out_payload_vaddr;
  wire                stage1Out_payload_tlb_hit;
  wire       [19:0]   stage1Out_payload_tlb_pageInfo_ppn;
  wire       [1:0]    stage1Out_payload_tlb_pageInfo_plv;
  wire       [1:0]    stage1Out_payload_tlb_pageInfo_mat;
  wire                stage1Out_payload_tlb_pageInfo_d;
  wire                stage1Out_payload_tlb_pageInfo_v;
  reg        [3:0]    stage1Out_payload_wayValid;
  reg        [3:0]    stage1Out_payload_wayDirty;
  wire                stage1Out_payload_isStoreTag;
  wire                stage1Out_payload_isIndexInvalidate;
  wire                stage1Out_payload_isHitInvalidate;
  wire                stage1Out_payload_checkTLBException;
  wire                stage1Out_payload_lsException;
  wire                stage2In_valid;
  wire                stage2In_ready;
  wire       [4:0]    stage2In_payload_robIdx;
  wire       [5:0]    stage2In_payload_prd;
  wire       [31:0]   stage2In_payload_branchResult_targetPC;
  wire                stage2In_payload_branchResult_branchResult;
  wire                stage2In_payload_branchResult_predictFail;
  wire                stage2In_payload_exceptionInfo_exception;
  wire       [5:0]    stage2In_payload_exceptionInfo_eCode;
  wire       [0:0]    stage2In_payload_exceptionInfo_eSubCode;
  wire       [31:0]   stage2In_payload_storeData;
  wire                stage2In_payload_lsCtrlBundle_load;
  wire                stage2In_payload_lsCtrlBundle_store;
  wire                stage2In_payload_lsCtrlBundle_signed;
  wire                stage2In_payload_lsCtrlBundle_ll;
  wire                stage2In_payload_lsCtrlBundle_sc;
  wire       [3:0]    stage2In_payload_lsCtrlBundle_lsMask;
  wire       [2:0]    stage2In_payload_lsCtrlBundle_size;
  wire                stage2In_payload_lsCtrlBundle_normalMemOp;
  wire       [31:0]   stage2In_payload_vaddr;
  wire                stage2In_payload_tlb_hit;
  wire       [19:0]   stage2In_payload_tlb_pageInfo_ppn;
  wire       [1:0]    stage2In_payload_tlb_pageInfo_plv;
  wire       [1:0]    stage2In_payload_tlb_pageInfo_mat;
  wire                stage2In_payload_tlb_pageInfo_d;
  wire                stage2In_payload_tlb_pageInfo_v;
  wire       [3:0]    stage2In_payload_wayValid;
  wire       [3:0]    stage2In_payload_wayDirty;
  wire                stage2In_payload_isStoreTag;
  wire                stage2In_payload_isIndexInvalidate;
  wire                stage2In_payload_isHitInvalidate;
  wire                stage2In_payload_checkTLBException;
  wire                stage2In_payload_lsException;
  reg                 stage1Out_thrown_valid;
  reg                 stage1Out_thrown_ready;
  wire       [4:0]    stage1Out_thrown_payload_robIdx;
  wire       [5:0]    stage1Out_thrown_payload_prd;
  wire       [31:0]   stage1Out_thrown_payload_branchResult_targetPC;
  wire                stage1Out_thrown_payload_branchResult_branchResult;
  wire                stage1Out_thrown_payload_branchResult_predictFail;
  wire                stage1Out_thrown_payload_exceptionInfo_exception;
  wire       [5:0]    stage1Out_thrown_payload_exceptionInfo_eCode;
  wire       [0:0]    stage1Out_thrown_payload_exceptionInfo_eSubCode;
  wire       [31:0]   stage1Out_thrown_payload_storeData;
  wire                stage1Out_thrown_payload_lsCtrlBundle_load;
  wire                stage1Out_thrown_payload_lsCtrlBundle_store;
  wire                stage1Out_thrown_payload_lsCtrlBundle_signed;
  wire                stage1Out_thrown_payload_lsCtrlBundle_ll;
  wire                stage1Out_thrown_payload_lsCtrlBundle_sc;
  wire       [3:0]    stage1Out_thrown_payload_lsCtrlBundle_lsMask;
  wire       [2:0]    stage1Out_thrown_payload_lsCtrlBundle_size;
  wire                stage1Out_thrown_payload_lsCtrlBundle_normalMemOp;
  wire       [31:0]   stage1Out_thrown_payload_vaddr;
  wire                stage1Out_thrown_payload_tlb_hit;
  wire       [19:0]   stage1Out_thrown_payload_tlb_pageInfo_ppn;
  wire       [1:0]    stage1Out_thrown_payload_tlb_pageInfo_plv;
  wire       [1:0]    stage1Out_thrown_payload_tlb_pageInfo_mat;
  wire                stage1Out_thrown_payload_tlb_pageInfo_d;
  wire                stage1Out_thrown_payload_tlb_pageInfo_v;
  wire       [3:0]    stage1Out_thrown_payload_wayValid;
  wire       [3:0]    stage1Out_thrown_payload_wayDirty;
  wire                stage1Out_thrown_payload_isStoreTag;
  wire                stage1Out_thrown_payload_isIndexInvalidate;
  wire                stage1Out_thrown_payload_isHitInvalidate;
  wire                stage1Out_thrown_payload_checkTLBException;
  wire                stage1Out_thrown_payload_lsException;
  wire                stage1Out_thrown_m2sPipe_valid;
  wire                stage1Out_thrown_m2sPipe_ready;
  wire       [4:0]    stage1Out_thrown_m2sPipe_payload_robIdx;
  wire       [5:0]    stage1Out_thrown_m2sPipe_payload_prd;
  wire       [31:0]   stage1Out_thrown_m2sPipe_payload_branchResult_targetPC;
  wire                stage1Out_thrown_m2sPipe_payload_branchResult_branchResult;
  wire                stage1Out_thrown_m2sPipe_payload_branchResult_predictFail;
  wire                stage1Out_thrown_m2sPipe_payload_exceptionInfo_exception;
  wire       [5:0]    stage1Out_thrown_m2sPipe_payload_exceptionInfo_eCode;
  wire       [0:0]    stage1Out_thrown_m2sPipe_payload_exceptionInfo_eSubCode;
  wire       [31:0]   stage1Out_thrown_m2sPipe_payload_storeData;
  wire                stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_load;
  wire                stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_store;
  wire                stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_signed;
  wire                stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_ll;
  wire                stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_sc;
  wire       [3:0]    stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_lsMask;
  wire       [2:0]    stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_size;
  wire                stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_normalMemOp;
  wire       [31:0]   stage1Out_thrown_m2sPipe_payload_vaddr;
  wire                stage1Out_thrown_m2sPipe_payload_tlb_hit;
  wire       [19:0]   stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_ppn;
  wire       [1:0]    stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_plv;
  wire       [1:0]    stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_mat;
  wire                stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_d;
  wire                stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_v;
  wire       [3:0]    stage1Out_thrown_m2sPipe_payload_wayValid;
  wire       [3:0]    stage1Out_thrown_m2sPipe_payload_wayDirty;
  wire                stage1Out_thrown_m2sPipe_payload_isStoreTag;
  wire                stage1Out_thrown_m2sPipe_payload_isIndexInvalidate;
  wire                stage1Out_thrown_m2sPipe_payload_isHitInvalidate;
  wire                stage1Out_thrown_m2sPipe_payload_checkTLBException;
  wire                stage1Out_thrown_m2sPipe_payload_lsException;
  reg                 stage1Out_thrown_rValid;
  reg        [4:0]    stage1Out_thrown_rData_robIdx;
  reg        [5:0]    stage1Out_thrown_rData_prd;
  reg        [31:0]   stage1Out_thrown_rData_branchResult_targetPC;
  reg                 stage1Out_thrown_rData_branchResult_branchResult;
  reg                 stage1Out_thrown_rData_branchResult_predictFail;
  reg                 stage1Out_thrown_rData_exceptionInfo_exception;
  reg        [5:0]    stage1Out_thrown_rData_exceptionInfo_eCode;
  reg        [0:0]    stage1Out_thrown_rData_exceptionInfo_eSubCode;
  reg        [31:0]   stage1Out_thrown_rData_storeData;
  reg                 stage1Out_thrown_rData_lsCtrlBundle_load;
  reg                 stage1Out_thrown_rData_lsCtrlBundle_store;
  reg                 stage1Out_thrown_rData_lsCtrlBundle_signed;
  reg                 stage1Out_thrown_rData_lsCtrlBundle_ll;
  reg                 stage1Out_thrown_rData_lsCtrlBundle_sc;
  reg        [3:0]    stage1Out_thrown_rData_lsCtrlBundle_lsMask;
  reg        [2:0]    stage1Out_thrown_rData_lsCtrlBundle_size;
  reg                 stage1Out_thrown_rData_lsCtrlBundle_normalMemOp;
  reg        [31:0]   stage1Out_thrown_rData_vaddr;
  reg                 stage1Out_thrown_rData_tlb_hit;
  reg        [19:0]   stage1Out_thrown_rData_tlb_pageInfo_ppn;
  reg        [1:0]    stage1Out_thrown_rData_tlb_pageInfo_plv;
  reg        [1:0]    stage1Out_thrown_rData_tlb_pageInfo_mat;
  reg                 stage1Out_thrown_rData_tlb_pageInfo_d;
  reg                 stage1Out_thrown_rData_tlb_pageInfo_v;
  reg        [3:0]    stage1Out_thrown_rData_wayValid;
  reg        [3:0]    stage1Out_thrown_rData_wayDirty;
  reg                 stage1Out_thrown_rData_isStoreTag;
  reg                 stage1Out_thrown_rData_isIndexInvalidate;
  reg                 stage1Out_thrown_rData_isHitInvalidate;
  reg                 stage1Out_thrown_rData_checkTLBException;
  reg                 stage1Out_thrown_rData_lsException;
  wire                when_Stream_l369;
  wire       [1:0]    preShiftSize;
  wire       [3:0]    switch_LSU_l94;
  reg        [25:0]   transferRAddrHi;
  reg        [3:0]    transferRAddrMid;
  reg        [1:0]    transferRAddrLo;
  wire       [31:0]   transferRAddr;
  reg        [25:0]   transferWAddrHi;
  reg        [3:0]    transferWAddrMid;
  reg        [1:0]    transferWAddrLo;
  wire       [31:0]   transferWAddr;
  reg                 transferUncached;
  reg                 transferCACOP;
  wire       [2:0]    transferWriteBufferIdx;
  reg        [31:0]   transferWData;
  reg        [3:0]    transferLSMask;
  reg        [3:0]    transferWaySelect;
  wire       [8:0]    portAddr0;
  reg        [31:0]   portRData0_0;
  reg        [31:0]   portRData0_1;
  reg        [31:0]   portRData0_2;
  reg        [31:0]   portRData0_3;
  wire       [31:0]   portRData0Raw_0;
  wire       [31:0]   portRData0Raw_1;
  wire       [31:0]   portRData0Raw_2;
  wire       [31:0]   portRData0Raw_3;
  wire       [31:0]   portWData0;
  wire       [3:0]    portWMask0;
  wire                portRen0_0;
  wire                portRen0_1;
  wire                portRen0_2;
  wire                portRen0_3;
  wire                portWen0_0;
  wire                portWen0_1;
  wire                portWen0_2;
  wire                portWen0_3;
  wire       [8:0]    portAddr1;
  wire       [31:0]   portRData1_0;
  wire       [31:0]   portRData1_1;
  wire       [31:0]   portRData1_2;
  wire       [31:0]   portRData1_3;
  wire       [31:0]   portWData1;
  wire       [3:0]    portWMask1;
  wire                portRen1_0;
  wire                portRen1_1;
  wire                portRen1_2;
  wire                portRen1_3;
  wire                portWen1_0;
  wire                portWen1_1;
  wire                portWen1_2;
  wire                portWen1_3;
  reg        [31:0]   portWData1Bypass_0;
  reg        [31:0]   portWData1Bypass_1;
  reg        [31:0]   portWData1Bypass_2;
  reg        [31:0]   portWData1Bypass_3;
  reg        [3:0]    portWMask1Bypass_0;
  reg        [3:0]    portWMask1Bypass_1;
  reg        [3:0]    portWMask1Bypass_2;
  reg        [3:0]    portWMask1Bypass_3;
  wire       [4:0]    missingEntry_robIdx;
  wire       [5:0]    missingEntry_prd;
  wire       [31:0]   missingEntry_branchResult_targetPC;
  wire                missingEntry_branchResult_branchResult;
  wire                missingEntry_branchResult_predictFail;
  wire                missingEntry_exceptionInfo_exception;
  wire       [5:0]    missingEntry_exceptionInfo_eCode;
  wire       [0:0]    missingEntry_exceptionInfo_eSubCode;
  wire                missingEntry_uncached;
  wire                missingEntry_load;
  wire                missingEntry_store;
  wire                missingEntry_signed;
  wire                missingEntry_ll;
  wire                missingEntry_sc;
  wire       [2:0]    missingEntry_writeBufferIdx;
  wire       [3:0]    missingEntry_waySelect;
  wire                missingEntry_writeBack;
  wire       [31:0]   missingEntry_storeData;
  wire       [3:0]    missingEntry_lsMask;
  wire       [2:0]    missingEntry_size;
  wire       [31:0]   missingEntry_vaddr;
  wire       [31:0]   missingEntry_paddr;
  wire       [31:0]   missingEntry_prevPaddr;
  wire                missingEntry_valid;
  wire       [4:0]    latestWrite_robIdx;
  wire       [3:0]    latestWrite_waySelect;
  wire       [31:0]   latestWrite_prevData;
  wire                latestWrite_prevDirty;
  wire       [8:0]    latestWrite_index;
  wire                latestWrite_miss;
  wire                latestWrite_valid;
  reg        [31:0]   mergedWrite;
  wire       [3:0]    _zz_portRen0_0;
  wire       [3:0]    _zz_portWen0_0;
  wire                _zz_portWen0_0_1;
  wire       [3:0]    _zz_portWen0_0_2;
  wire                _zz_portRen1_0;
  wire       [3:0]    _zz_portRen1_0_1;
  wire                _zz_portWen1_1;
  wire                _zz_portWen1_2;
  wire                _zz_portWen1_3;
  wire                _zz_portWen1_0;
  wire       [3:0]    _zz_portWen1_0_1;
  wire                _zz_portWen1_1_1;
  wire                _zz_portWen1_2_1;
  wire                _zz_portWen1_3_1;
  wire                _zz_portWen1_0_2;
  wire       [3:0]    _zz_portWen1_0_3;
  wire       [3:0]    _zz_portWen1_0_4;
  wire                _zz_portWen1_0_5;
  wire       [3:0]    _zz_portWen1_0_6;
  wire                when_LSU_l174;
  wire                when_LSU_l174_1;
  wire                when_LSU_l174_2;
  wire                when_LSU_l174_3;
  wire                stage1Out_fire;
  wire                _zz_exceptionInfo_exception;
  wire                hasException;
  reg                 axiLoad;
  reg                 axiFinish;
  wire                noStructuralHazard;
  wire                when_LSU_l203;
  wire                when_LSU_l213;
  wire                when_LSU_l217;
  wire                when_LSU_l221;
  wire                scMatchHit;
  wire                scMatchAXI;
  wire       [31:0]   scResHit;
  wire       [31:0]   scResAXI;
  reg        [7:0]    writeBufferRetireMask;
  reg        [4:0]    writeBuffer_0_robIdx;
  reg        [3:0]    writeBuffer_0_waySelect;
  reg        [31:0]   writeBuffer_0_prevData;
  reg                 writeBuffer_0_prevDirty;
  reg        [8:0]    writeBuffer_0_index;
  reg                 writeBuffer_0_miss;
  reg                 writeBuffer_0_valid;
  reg        [4:0]    writeBuffer_1_robIdx;
  reg        [3:0]    writeBuffer_1_waySelect;
  reg        [31:0]   writeBuffer_1_prevData;
  reg                 writeBuffer_1_prevDirty;
  reg        [8:0]    writeBuffer_1_index;
  reg                 writeBuffer_1_miss;
  reg                 writeBuffer_1_valid;
  reg        [4:0]    writeBuffer_2_robIdx;
  reg        [3:0]    writeBuffer_2_waySelect;
  reg        [31:0]   writeBuffer_2_prevData;
  reg                 writeBuffer_2_prevDirty;
  reg        [8:0]    writeBuffer_2_index;
  reg                 writeBuffer_2_miss;
  reg                 writeBuffer_2_valid;
  reg        [4:0]    writeBuffer_3_robIdx;
  reg        [3:0]    writeBuffer_3_waySelect;
  reg        [31:0]   writeBuffer_3_prevData;
  reg                 writeBuffer_3_prevDirty;
  reg        [8:0]    writeBuffer_3_index;
  reg                 writeBuffer_3_miss;
  reg                 writeBuffer_3_valid;
  reg        [4:0]    writeBuffer_4_robIdx;
  reg        [3:0]    writeBuffer_4_waySelect;
  reg        [31:0]   writeBuffer_4_prevData;
  reg                 writeBuffer_4_prevDirty;
  reg        [8:0]    writeBuffer_4_index;
  reg                 writeBuffer_4_miss;
  reg                 writeBuffer_4_valid;
  reg        [4:0]    writeBuffer_5_robIdx;
  reg        [3:0]    writeBuffer_5_waySelect;
  reg        [31:0]   writeBuffer_5_prevData;
  reg                 writeBuffer_5_prevDirty;
  reg        [8:0]    writeBuffer_5_index;
  reg                 writeBuffer_5_miss;
  reg                 writeBuffer_5_valid;
  reg        [4:0]    writeBuffer_6_robIdx;
  reg        [3:0]    writeBuffer_6_waySelect;
  reg        [31:0]   writeBuffer_6_prevData;
  reg                 writeBuffer_6_prevDirty;
  reg        [8:0]    writeBuffer_6_index;
  reg                 writeBuffer_6_miss;
  reg                 writeBuffer_6_valid;
  reg        [4:0]    writeBuffer_7_robIdx;
  reg        [3:0]    writeBuffer_7_waySelect;
  reg        [31:0]   writeBuffer_7_prevData;
  reg                 writeBuffer_7_prevDirty;
  reg        [8:0]    writeBuffer_7_index;
  reg                 writeBuffer_7_miss;
  reg                 writeBuffer_7_valid;
  reg        [2:0]    writeBufferHead;
  reg        [2:0]    writeBufferTail;
  wire       [3:0]    _zz_writeBufferHeadNext;
  wire       [3:0]    _zz_writeBufferHeadNext_1;
  wire       [3:0]    _zz_writeBufferHeadNext_2;
  wire       [3:0]    _zz_writeBufferHeadNext_3;
  wire       [3:0]    _zz_writeBufferHeadNext_4;
  wire       [3:0]    _zz_writeBufferHeadNext_5;
  wire       [3:0]    _zz_writeBufferHeadNext_6;
  wire       [3:0]    _zz_writeBufferHeadNext_7;
  wire       [2:0]    writeBufferHeadNext;
  wire                _zz_writeBufferAvail;
  wire       [7:0]    _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  reg        [1:0]    _zz_writeBufferRetireMask;
  reg        [1:0]    _zz_writeBufferRetireMask_1;
  reg        [1:0]    _zz_writeBufferRetireMask_2;
  reg        [1:0]    _zz_writeBufferRetireMask_3;
  reg        [1:0]    _zz_writeBufferRetireMask_4;
  reg        [1:0]    _zz_writeBufferRetireMask_5;
  reg        [1:0]    _zz_writeBufferRetireMask_6;
  reg        [1:0]    _zz_writeBufferRetireMask_7;
  wire                when_LSU_l267;
  wire       [3:0]    _zz_writeBuffer_0_waySelect;
  wire                _zz_io_output_payload_data;
  wire                _zz_io_output_payload_data_1;
  wire       [1:0]    _zz_io_output_payload_data_2;
  wire       [31:0]   _zz_writeBuffer_0_prevData;
  wire                _zz_missBuffer_0_writeBack;
  wire                _zz_missBuffer_0_writeBack_1;
  wire                _zz_missBuffer_0_writeBack_2;
  wire                _zz_missBuffer_0_writeBack_3;
  wire                _zz_writeBuffer_0_prevDirty;
  wire       [8:0]    _zz_writeBuffer_0_index;
  wire       [7:0]    _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  reg        [4:0]    missBuffer_0_robIdx;
  reg        [5:0]    missBuffer_0_prd;
  reg        [31:0]   missBuffer_0_branchResult_targetPC;
  reg                 missBuffer_0_branchResult_branchResult;
  reg                 missBuffer_0_branchResult_predictFail;
  reg                 missBuffer_0_exceptionInfo_exception;
  reg        [5:0]    missBuffer_0_exceptionInfo_eCode;
  reg        [0:0]    missBuffer_0_exceptionInfo_eSubCode;
  reg                 missBuffer_0_uncached;
  reg                 missBuffer_0_load;
  reg                 missBuffer_0_store;
  reg                 missBuffer_0_signed;
  reg                 missBuffer_0_ll;
  reg                 missBuffer_0_sc;
  reg        [2:0]    missBuffer_0_writeBufferIdx;
  reg        [3:0]    missBuffer_0_waySelect;
  reg                 missBuffer_0_writeBack;
  reg        [31:0]   missBuffer_0_storeData;
  reg        [3:0]    missBuffer_0_lsMask;
  reg        [2:0]    missBuffer_0_size;
  reg        [31:0]   missBuffer_0_vaddr;
  reg        [31:0]   missBuffer_0_paddr;
  reg        [31:0]   missBuffer_0_prevPaddr;
  reg                 missBuffer_0_valid;
  wire                _zz_19;
  wire                when_LSU_l292;
  wire                _zz_missBuffer_0_writeBack_4;
  wire                _zz_missBuffer_0_writeBack_5;
  wire                _zz_missBuffer_0_writeBack_6;
  wire       [1:0]    _zz_missBuffer_0_writeBack_7;
  reg        [1:0]    sameBlockMask;
  wire                sameBlock;
  reg                 lruBit_0_0;
  reg                 lruBit_0_1;
  reg                 lruBit_0_2;
  reg                 lruBit_1_0;
  reg                 lruBit_1_1;
  reg                 lruBit_1_2;
  reg                 lruBit_2_0;
  reg                 lruBit_2_1;
  reg                 lruBit_2_2;
  reg                 lruBit_3_0;
  reg                 lruBit_3_1;
  reg                 lruBit_3_2;
  reg                 lruBit_4_0;
  reg                 lruBit_4_1;
  reg                 lruBit_4_2;
  reg                 lruBit_5_0;
  reg                 lruBit_5_1;
  reg                 lruBit_5_2;
  reg                 lruBit_6_0;
  reg                 lruBit_6_1;
  reg                 lruBit_6_2;
  reg                 lruBit_7_0;
  reg                 lruBit_7_1;
  reg                 lruBit_7_2;
  reg                 lruBit_8_0;
  reg                 lruBit_8_1;
  reg                 lruBit_8_2;
  reg                 lruBit_9_0;
  reg                 lruBit_9_1;
  reg                 lruBit_9_2;
  reg                 lruBit_10_0;
  reg                 lruBit_10_1;
  reg                 lruBit_10_2;
  reg                 lruBit_11_0;
  reg                 lruBit_11_1;
  reg                 lruBit_11_2;
  reg                 lruBit_12_0;
  reg                 lruBit_12_1;
  reg                 lruBit_12_2;
  reg                 lruBit_13_0;
  reg                 lruBit_13_1;
  reg                 lruBit_13_2;
  reg                 lruBit_14_0;
  reg                 lruBit_14_1;
  reg                 lruBit_14_2;
  reg                 lruBit_15_0;
  reg                 lruBit_15_1;
  reg                 lruBit_15_2;
  reg                 lruBit_16_0;
  reg                 lruBit_16_1;
  reg                 lruBit_16_2;
  reg                 lruBit_17_0;
  reg                 lruBit_17_1;
  reg                 lruBit_17_2;
  reg                 lruBit_18_0;
  reg                 lruBit_18_1;
  reg                 lruBit_18_2;
  reg                 lruBit_19_0;
  reg                 lruBit_19_1;
  reg                 lruBit_19_2;
  reg                 lruBit_20_0;
  reg                 lruBit_20_1;
  reg                 lruBit_20_2;
  reg                 lruBit_21_0;
  reg                 lruBit_21_1;
  reg                 lruBit_21_2;
  reg                 lruBit_22_0;
  reg                 lruBit_22_1;
  reg                 lruBit_22_2;
  reg                 lruBit_23_0;
  reg                 lruBit_23_1;
  reg                 lruBit_23_2;
  reg                 lruBit_24_0;
  reg                 lruBit_24_1;
  reg                 lruBit_24_2;
  reg                 lruBit_25_0;
  reg                 lruBit_25_1;
  reg                 lruBit_25_2;
  reg                 lruBit_26_0;
  reg                 lruBit_26_1;
  reg                 lruBit_26_2;
  reg                 lruBit_27_0;
  reg                 lruBit_27_1;
  reg                 lruBit_27_2;
  reg                 lruBit_28_0;
  reg                 lruBit_28_1;
  reg                 lruBit_28_2;
  reg                 lruBit_29_0;
  reg                 lruBit_29_1;
  reg                 lruBit_29_2;
  reg                 lruBit_30_0;
  reg                 lruBit_30_1;
  reg                 lruBit_30_2;
  reg                 lruBit_31_0;
  reg                 lruBit_31_1;
  reg                 lruBit_31_2;
  wire                io_output_fire;
  wire                when_LSU_l335;
  wire       [31:0]   _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_lruBit_0_0;
  wire                _zz_lruBit_0_1;
  wire                _zz_lruBit_0_2;
  wire                dirtyUpdate;
  wire                when_LSU_l341;
  wire       [31:0]   _zz_53;
  wire                when_LSU_l341_1;
  wire       [31:0]   _zz_54;
  wire                when_LSU_l341_2;
  wire       [31:0]   _zz_55;
  wire                when_LSU_l341_3;
  wire       [31:0]   _zz_56;
  wire                when_LSU_l348;
  wire       [31:0]   _zz_57;
  wire                when_LSU_l348_1;
  wire       [31:0]   _zz_58;
  wire                when_LSU_l348_2;
  wire       [31:0]   _zz_59;
  wire                when_LSU_l348_3;
  wire       [31:0]   _zz_60;
  wire                when_LSU_l357;
  wire                _zz_io_axi_wdata;
  wire                _zz_io_axi_wdata_1;
  wire       [0:0]    missBufferAllowMask;
  wire       [0:0]    missBufferPreAllowMask;
  reg        [1:0]    _zz_missBufferAllowMask;
  reg        [7:0]    _zz_missBufferPreAllowMask;
  wire       [31:0]   cacopPAddr;
  wire                axiCtrl_wantExit;
  reg                 axiCtrl_wantStart;
  wire                axiCtrl_wantKill;
  wire                rollbackCtrl_wantExit;
  reg                 rollbackCtrl_wantStart;
  wire                rollbackCtrl_wantKill;
  reg        [1:0]    _zz_wayToReplace;
  reg        [1:0]    _zz_wayToReplace_1;
  reg        [1:0]    _zz_wayToReplace_2;
  reg        [1:0]    _zz_wayToReplace_3;
  reg        [31:0]   dataShuffle_0;
  reg        [31:0]   dataShuffle_1;
  reg        [31:0]   dataShuffle_2;
  reg        [31:0]   dataShuffle_3;
  reg        [31:0]   axiShuffle;
  wire       [31:0]   _zz_dataShuffle_0;
  wire                _zz_dataShuffle_0_1;
  wire                _zz_dataShuffle_0_2;
  wire       [31:0]   _zz_dataShuffle_1;
  wire                _zz_dataShuffle_1_1;
  wire                _zz_dataShuffle_1_2;
  wire       [31:0]   _zz_dataShuffle_2;
  wire                _zz_dataShuffle_2_1;
  wire                _zz_dataShuffle_2_2;
  wire       [31:0]   _zz_dataShuffle_3;
  wire                _zz_dataShuffle_3_1;
  wire                _zz_dataShuffle_3_2;
  wire       [31:0]   axiShiftedData;
  wire                _zz_axiShuffle;
  wire                _zz_axiShuffle_1;
  wire       [4:0]    cacopIdx;
  wire       [3:0]    cacopWay;
  reg                 cacopWriteBack;
  wire                cacopSetInvalid;
  wire                when_LSU_l661;
  wire                when_LSU_l663;
  wire       [31:0]   _zz_61;
  wire                when_LSU_l663_1;
  wire       [31:0]   _zz_62;
  wire                when_LSU_l663_2;
  wire       [31:0]   _zz_63;
  wire                when_LSU_l663_3;
  wire       [31:0]   _zz_64;
  wire                specialOpBufferWrite;
  reg        [2:0]    axiCtrl_stateReg;
  reg        [2:0]    axiCtrl_stateNext;
  wire                when_LSU_l436;
  wire                when_LSU_l447;
  wire                when_LSU_l453;
  wire                when_LSU_l471;
  wire                when_LSU_l473;
  wire       [31:0]   _zz_65;
  wire       [31:0]   _zz_66;
  wire                when_LSU_l473_1;
  wire       [31:0]   _zz_67;
  wire       [31:0]   _zz_68;
  wire                when_LSU_l473_2;
  wire       [31:0]   _zz_69;
  wire       [31:0]   _zz_70;
  wire                when_LSU_l473_3;
  wire       [31:0]   _zz_71;
  wire       [31:0]   _zz_72;
  wire                when_LSU_l480;
  wire                when_LSU_l481;
  wire                when_LSU_l496;
  wire                when_LSU_l510;
  wire                when_LSU_l527;
  wire                when_LSU_l539;
  reg        [1:0]    rollbackCtrl_stateReg;
  reg        [1:0]    rollbackCtrl_stateNext;
  wire                when_LSU_l564;
  wire                when_LSU_l567;
  wire                when_LSU_l575;
  `ifndef SYNTHESIS
  reg [55:0] io_input_payload_uop_lsuOp_string;
  reg [55:0] io_specialOpBufferUpdate_payload_uop_lsuOp_string;
  reg [71:0] axiCtrl_stateReg_string;
  reg [71:0] axiCtrl_stateNext_string;
  reg [63:0] rollbackCtrl_stateReg_string;
  reg [63:0] rollbackCtrl_stateNext_string;
  `endif


  assign _zz_stage1Out_payload_storeData = (io_input_payload_src3 <<< preShiftSize);
  assign _zz_stage1Out_payload_lsCtrlBundle_size = 1'b1;
  assign _zz_stage1Out_payload_lsCtrlBundle_size_1 = 2'b10;
  assign _zz_stage1Out_payload_lsCtrlBundle_size_2 = 2'b10;
  assign _zz_stage1Out_payload_checkTLBException_1 = 2'b10;
  assign _zz_stage1Out_payload_checkTLBException = {3'd0, _zz_stage1Out_payload_checkTLBException_1};
  assign _zz_portAddr0 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : address);
  assign _zz_portAddr1 = transferRAddr;
  assign _zz_portAddr1_1 = transferWAddr;
  assign _zz_stage1Out_payload_wayValid_2 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_stage1Out_payload_wayDirty_2 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_hit_1 = 1'b1;
  assign _zz_hit = {1'd0, _zz_hit_1};
  assign _zz_stage1Out_payload_wayValid_5 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_stage1Out_payload_wayDirty_5 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_hit_3 = 1'b1;
  assign _zz_hit_2 = {1'd0, _zz_hit_3};
  assign _zz_stage1Out_payload_wayValid_8 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_stage1Out_payload_wayDirty_8 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_hit_5 = 1'b1;
  assign _zz_hit_4 = {1'd0, _zz_hit_5};
  assign _zz_stage1Out_payload_wayValid_11 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_stage1Out_payload_wayDirty_11 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_hit_7 = 1'b1;
  assign _zz_hit_6 = {1'd0, _zz_hit_7};
  assign _zz_exceptionInfo1_eCode = 4'b1001;
  assign _zz_exceptionInfo1_eCode_1 = 4'b1001;
  assign _zz_exceptionInfo2_eCode_1 = 1'b1;
  assign _zz_exceptionInfo2_eCode = {5'd0, _zz_exceptionInfo2_eCode_1};
  assign _zz_exceptionInfo2_eCode_3 = 2'b10;
  assign _zz_exceptionInfo2_eCode_2 = {4'd0, _zz_exceptionInfo2_eCode_3};
  assign _zz_exceptionInfo2_eCode_4 = 3'b111;
  assign _zz_exceptionInfo2_eCode_5 = 3'b100;
  assign _zz_exceptionInfo2_eCode_6 = 3'b111;
  assign _zz_writeBufferHeadNext_9 = (_zz_writeBufferHeadNext_10 + _zz_writeBufferHeadNext_15);
  assign _zz_writeBufferHeadNext_8 = _zz_writeBufferHeadNext_9[2:0];
  assign _zz_writeBufferHeadNext_10 = (_zz_writeBufferHeadNext_11 + _zz_writeBufferHeadNext_13);
  assign _zz_writeBufferHeadNext_17 = {writeBufferRetireMask[7],writeBufferRetireMask[6]};
  assign _zz_writeBufferHeadNext_16 = {1'd0, _zz_writeBufferHeadNext_17};
  assign _zz_writeBufferAppend_1 = 1'b1;
  assign _zz_writeBufferAppend = {1'd0, _zz_writeBufferAppend_1};
  assign _zz__zz_19 = 1'b1;
  assign _zz_when_LSU_l335_1 = 1'b1;
  assign _zz_when_LSU_l335 = {1'd0, _zz_when_LSU_l335_1};
  assign _zz_dirtyUpdate_1 = 1'b1;
  assign _zz_dirtyUpdate = {1'd0, _zz_dirtyUpdate_1};
  assign _zz__zz_53 = transferRAddr;
  assign _zz__zz_54 = transferRAddr;
  assign _zz__zz_55 = transferRAddr;
  assign _zz__zz_56 = transferRAddr;
  assign _zz_when_LSU_l357 = transferRAddr;
  assign _zz_when_LSU_l357_1 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_io_axi_arid = 1'b1;
  assign _zz_io_axi_arlen_1 = 4'b1111;
  assign _zz_io_axi_arlen = {4'd0, _zz_io_axi_arlen_1};
  assign _zz_io_axi_arsize_1 = 2'b10;
  assign _zz_io_axi_arsize = {1'd0, _zz_io_axi_arsize_1};
  assign _zz_io_axi_awid = 1'b1;
  assign _zz_io_axi_awlen = 4'b1111;
  assign _zz_io_axi_awsize_1 = 2'b10;
  assign _zz_io_axi_awsize = {1'd0, _zz_io_axi_awsize_1};
  assign _zz_io_axi_awburst = 1'b1;
  assign _zz_io_axi_wid = 1'b1;
  assign _zz__zz_missBufferAllowMask = {io_retireComm_allowRetire_1,io_retireComm_allowRetire_0};
  assign _zz__zz_missBufferPreAllowMask_1 = missBuffer_0_vaddr[10 : 6];
  assign _zz__zz_missBufferPreAllowMask = {4'd0, _zz__zz_missBufferPreAllowMask_1};
  assign _zz__zz_missBufferPreAllowMask_3 = missBuffer_0_vaddr[10 : 6];
  assign _zz__zz_missBufferPreAllowMask_2 = {4'd0, _zz__zz_missBufferPreAllowMask_3};
  assign _zz__zz_missBufferPreAllowMask_5 = missBuffer_0_vaddr[10 : 6];
  assign _zz__zz_missBufferPreAllowMask_4 = {4'd0, _zz__zz_missBufferPreAllowMask_5};
  assign _zz__zz_missBufferPreAllowMask_7 = missBuffer_0_vaddr[10 : 6];
  assign _zz__zz_missBufferPreAllowMask_6 = {4'd0, _zz__zz_missBufferPreAllowMask_7};
  assign _zz__zz_missBufferPreAllowMask_9 = missBuffer_0_vaddr[10 : 6];
  assign _zz__zz_missBufferPreAllowMask_8 = {4'd0, _zz__zz_missBufferPreAllowMask_9};
  assign _zz__zz_missBufferPreAllowMask_11 = missBuffer_0_vaddr[10 : 6];
  assign _zz__zz_missBufferPreAllowMask_10 = {4'd0, _zz__zz_missBufferPreAllowMask_11};
  assign _zz__zz_missBufferPreAllowMask_13 = missBuffer_0_vaddr[10 : 6];
  assign _zz__zz_missBufferPreAllowMask_12 = {4'd0, _zz__zz_missBufferPreAllowMask_13};
  assign _zz__zz_missBufferPreAllowMask_15 = missBuffer_0_vaddr[10 : 6];
  assign _zz__zz_missBufferPreAllowMask_14 = {4'd0, _zz__zz_missBufferPreAllowMask_15};
  assign _zz_cacopWay = (4'b0001 <<< stage2In_payload_vaddr[1 : 0]);
  assign _zz__zz_65 = transferRAddr;
  assign _zz__zz_66 = transferRAddr;
  assign _zz__zz_67 = transferRAddr;
  assign _zz__zz_68 = transferRAddr;
  assign _zz__zz_69 = transferRAddr;
  assign _zz__zz_70 = transferRAddr;
  assign _zz__zz_71 = transferRAddr;
  assign _zz__zz_72 = transferRAddr;
  assign _zz_transferRAddrMid = (transferRAddrMid + 4'b0001);
  assign _zz_transferRAddrMid_1 = (transferRAddrMid + 4'b0001);
  assign _zz_transferWAddrMid = (transferWAddrMid + 4'b0001);
  assign _zz_wr_addr = transferRAddr;
  assign _zz_wr_data = transferRAddr;
  assign _zz_rd_addr = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_wr_addr_1 = transferRAddr;
  assign _zz_wr_data_1 = transferRAddr;
  assign _zz_rd_addr_1 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_wr_addr_2 = transferRAddr;
  assign _zz_wr_data_2 = transferRAddr;
  assign _zz_rd_addr_2 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_wr_addr_3 = transferRAddr;
  assign _zz_wr_data_3 = transferRAddr;
  assign _zz_rd_addr_3 = (cacopEn ? io_ctrl_cacopVA : address);
  assign _zz_stage1Out_payload_wayValid_1 = _zz_stage1Out_payload_wayValid_2[10 : 6];
  assign _zz_stage1Out_payload_wayDirty_1 = _zz_stage1Out_payload_wayDirty_2[10 : 6];
  assign _zz_stage1Out_payload_wayValid_4 = _zz_stage1Out_payload_wayValid_5[10 : 6];
  assign _zz_stage1Out_payload_wayDirty_4 = _zz_stage1Out_payload_wayDirty_5[10 : 6];
  assign _zz_stage1Out_payload_wayValid_7 = _zz_stage1Out_payload_wayValid_8[10 : 6];
  assign _zz_stage1Out_payload_wayDirty_7 = _zz_stage1Out_payload_wayDirty_8[10 : 6];
  assign _zz_stage1Out_payload_wayValid_10 = _zz_stage1Out_payload_wayValid_11[10 : 6];
  assign _zz_stage1Out_payload_wayDirty_10 = _zz_stage1Out_payload_wayDirty_11[10 : 6];
  assign _zz_writeBufferHeadNext_12 = {writeBufferRetireMask[2],{writeBufferRetireMask[1],writeBufferRetireMask[0]}};
  assign _zz_writeBufferHeadNext_14 = {writeBufferRetireMask[5],{writeBufferRetireMask[4],writeBufferRetireMask[3]}};
  assign _zz_io_axi_wdata_3 = {_zz_io_axi_wdata_1,_zz_io_axi_wdata};
  assign _zz_cacopPAddr_1 = stage2In_payload_vaddr[1 : 0];
  assign _zz__zz_wayToReplace_1 = stage2In_payload_vaddr[10 : 6];
  assign _zz__zz_wayToReplace_3 = stage2In_payload_vaddr[10 : 6];
  assign _zz__zz_wayToReplace_1_2 = stage2In_payload_vaddr[10 : 6];
  assign _zz__zz_wayToReplace_1_4 = stage2In_payload_vaddr[10 : 6];
  assign _zz__zz_wayToReplace_2_2 = stage2In_payload_vaddr[10 : 6];
  assign _zz__zz_wayToReplace_2_4 = stage2In_payload_vaddr[10 : 6];
  assign _zz__zz_wayToReplace_3_2 = stage2In_payload_vaddr[10 : 6];
  assign _zz__zz_wayToReplace_3_4 = stage2In_payload_vaddr[10 : 6];
  assign _zz_dataShuffle_0_3 = _zz_dataShuffle_0_1;
  assign _zz_dataShuffle_0_4 = {_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,_zz_dataShuffle_0_1}}}}}}}}}}}}};
  assign _zz_dataShuffle_0_5 = _zz_dataShuffle_0_2;
  assign _zz_dataShuffle_0_6 = {_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,_zz_dataShuffle_0_2}}}}};
  assign _zz_dataShuffle_1_3 = _zz_dataShuffle_1_1;
  assign _zz_dataShuffle_1_4 = {_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,_zz_dataShuffle_1_1}}}}}}}}}}}}};
  assign _zz_dataShuffle_1_5 = _zz_dataShuffle_1_2;
  assign _zz_dataShuffle_1_6 = {_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,_zz_dataShuffle_1_2}}}}};
  assign _zz_dataShuffle_2_3 = _zz_dataShuffle_2_1;
  assign _zz_dataShuffle_2_4 = {_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,_zz_dataShuffle_2_1}}}}}}}}}}}}};
  assign _zz_dataShuffle_2_5 = _zz_dataShuffle_2_2;
  assign _zz_dataShuffle_2_6 = {_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,_zz_dataShuffle_2_2}}}}};
  assign _zz_dataShuffle_3_3 = _zz_dataShuffle_3_1;
  assign _zz_dataShuffle_3_4 = {_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,_zz_dataShuffle_3_1}}}}}}}}}}}}};
  assign _zz_dataShuffle_3_5 = _zz_dataShuffle_3_2;
  assign _zz_dataShuffle_3_6 = {_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,_zz_dataShuffle_3_2}}}}};
  assign _zz_axiShuffle_2 = _zz_axiShuffle;
  assign _zz_axiShuffle_3 = {_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,_zz_axiShuffle}}}}}}}}}}}}};
  assign _zz_axiShuffle_4 = _zz_axiShuffle_1;
  assign _zz_axiShuffle_5 = {_zz_axiShuffle_1,{_zz_axiShuffle_1,{_zz_axiShuffle_1,{_zz_axiShuffle_1,{_zz_axiShuffle_1,_zz_axiShuffle_1}}}}};
  Ram_2wrs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .portA_readUnderWrite("dontCare"),
    .portA_duringWrite("dontCare"),
    .portA_addressWidth(9),
    .portA_dataWidth(32),
    .portA_maskWidth(4),
    .portA_maskEnable(1'b1),
    .portB_readUnderWrite("dontCare"),
    .portB_duringWrite("dontCare"),
    .portB_addressWidth(9),
    .portB_dataWidth(32),
    .portB_maskWidth(4),
    .portB_maskEnable(1'b1)
  ) data_0 (
    .portA_clk    (aclk                     ), //i
    .portA_en     (data_0_portA_en          ), //i
    .portA_wr     (portWen0_0               ), //i
    .portA_mask   (portWMask0[3:0]          ), //i
    .portA_addr   (portAddr0[8:0]           ), //i
    .portA_wrData (portWData0[31:0]         ), //i
    .portA_rdData (data_0_portA_rdData[31:0]), //o
    .portB_clk    (aclk                     ), //i
    .portB_en     (data_0_portB_en          ), //i
    .portB_wr     (portWen1_0               ), //i
    .portB_mask   (portWMask1[3:0]          ), //i
    .portB_addr   (portAddr1[8:0]           ), //i
    .portB_wrData (portWData1[31:0]         ), //i
    .portB_rdData (data_0_portB_rdData[31:0])  //o
  );
  Ram_2wrs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .portA_readUnderWrite("dontCare"),
    .portA_duringWrite("dontCare"),
    .portA_addressWidth(9),
    .portA_dataWidth(32),
    .portA_maskWidth(4),
    .portA_maskEnable(1'b1),
    .portB_readUnderWrite("dontCare"),
    .portB_duringWrite("dontCare"),
    .portB_addressWidth(9),
    .portB_dataWidth(32),
    .portB_maskWidth(4),
    .portB_maskEnable(1'b1)
  ) data_1 (
    .portA_clk    (aclk                     ), //i
    .portA_en     (data_1_portA_en          ), //i
    .portA_wr     (portWen0_1               ), //i
    .portA_mask   (portWMask0[3:0]          ), //i
    .portA_addr   (portAddr0[8:0]           ), //i
    .portA_wrData (portWData0[31:0]         ), //i
    .portA_rdData (data_1_portA_rdData[31:0]), //o
    .portB_clk    (aclk                     ), //i
    .portB_en     (data_1_portB_en          ), //i
    .portB_wr     (portWen1_1               ), //i
    .portB_mask   (portWMask1[3:0]          ), //i
    .portB_addr   (portAddr1[8:0]           ), //i
    .portB_wrData (portWData1[31:0]         ), //i
    .portB_rdData (data_1_portB_rdData[31:0])  //o
  );
  Ram_2wrs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .portA_readUnderWrite("dontCare"),
    .portA_duringWrite("dontCare"),
    .portA_addressWidth(9),
    .portA_dataWidth(32),
    .portA_maskWidth(4),
    .portA_maskEnable(1'b1),
    .portB_readUnderWrite("dontCare"),
    .portB_duringWrite("dontCare"),
    .portB_addressWidth(9),
    .portB_dataWidth(32),
    .portB_maskWidth(4),
    .portB_maskEnable(1'b1)
  ) data_2 (
    .portA_clk    (aclk                     ), //i
    .portA_en     (data_2_portA_en          ), //i
    .portA_wr     (portWen0_2               ), //i
    .portA_mask   (portWMask0[3:0]          ), //i
    .portA_addr   (portAddr0[8:0]           ), //i
    .portA_wrData (portWData0[31:0]         ), //i
    .portA_rdData (data_2_portA_rdData[31:0]), //o
    .portB_clk    (aclk                     ), //i
    .portB_en     (data_2_portB_en          ), //i
    .portB_wr     (portWen1_2               ), //i
    .portB_mask   (portWMask1[3:0]          ), //i
    .portB_addr   (portAddr1[8:0]           ), //i
    .portB_wrData (portWData1[31:0]         ), //i
    .portB_rdData (data_2_portB_rdData[31:0])  //o
  );
  Ram_2wrs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .portA_readUnderWrite("dontCare"),
    .portA_duringWrite("dontCare"),
    .portA_addressWidth(9),
    .portA_dataWidth(32),
    .portA_maskWidth(4),
    .portA_maskEnable(1'b1),
    .portB_readUnderWrite("dontCare"),
    .portB_duringWrite("dontCare"),
    .portB_addressWidth(9),
    .portB_dataWidth(32),
    .portB_maskWidth(4),
    .portB_maskEnable(1'b1)
  ) data_3 (
    .portA_clk    (aclk                     ), //i
    .portA_en     (data_3_portA_en          ), //i
    .portA_wr     (portWen0_3               ), //i
    .portA_mask   (portWMask0[3:0]          ), //i
    .portA_addr   (portAddr0[8:0]           ), //i
    .portA_wrData (portWData0[31:0]         ), //i
    .portA_rdData (data_3_portA_rdData[31:0]), //o
    .portB_clk    (aclk                     ), //i
    .portB_en     (data_3_portB_en          ), //i
    .portB_wr     (portWen1_3               ), //i
    .portB_mask   (portWMask1[3:0]          ), //i
    .portB_addr   (portAddr1[8:0]           ), //i
    .portB_wrData (portWData1[31:0]         ), //i
    .portB_rdData (data_3_portB_rdData[31:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_0 (
    .wr_clk  (aclk               ), //i
    .wr_en   (tag_0_wr_en        ), //i
    .wr_mask (tag_0_wr_mask      ), //i
    .wr_addr (tag_0_wr_addr[4:0] ), //i
    .wr_data (tag_0_wr_data[20:0]), //i
    .rd_clk  (aclk               ), //i
    .rd_en   (tag_0_rd_en        ), //i
    .rd_addr (tag_0_rd_addr[4:0] ), //i
    .rd_data (tag_0_rd_data[20:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_1 (
    .wr_clk  (aclk               ), //i
    .wr_en   (tag_1_wr_en        ), //i
    .wr_mask (tag_1_wr_mask      ), //i
    .wr_addr (tag_1_wr_addr[4:0] ), //i
    .wr_data (tag_1_wr_data[20:0]), //i
    .rd_clk  (aclk               ), //i
    .rd_en   (tag_1_rd_en        ), //i
    .rd_addr (tag_1_rd_addr[4:0] ), //i
    .rd_data (tag_1_rd_data[20:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_2 (
    .wr_clk  (aclk               ), //i
    .wr_en   (tag_2_wr_en        ), //i
    .wr_mask (tag_2_wr_mask      ), //i
    .wr_addr (tag_2_wr_addr[4:0] ), //i
    .wr_data (tag_2_wr_data[20:0]), //i
    .rd_clk  (aclk               ), //i
    .rd_en   (tag_2_rd_en        ), //i
    .rd_addr (tag_2_rd_addr[4:0] ), //i
    .rd_data (tag_2_rd_data[20:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_3 (
    .wr_clk  (aclk               ), //i
    .wr_en   (tag_3_wr_en        ), //i
    .wr_mask (tag_3_wr_mask      ), //i
    .wr_addr (tag_3_wr_addr[4:0] ), //i
    .wr_data (tag_3_wr_data[20:0]), //i
    .rd_clk  (aclk               ), //i
    .rd_en   (tag_3_rd_en        ), //i
    .rd_addr (tag_3_rd_addr[4:0] ), //i
    .rd_data (tag_3_rd_data[20:0])  //o
  );
  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_1)
      5'b00000 : _zz_stage1Out_payload_wayValid = valid_0_0;
      5'b00001 : _zz_stage1Out_payload_wayValid = valid_0_1;
      5'b00010 : _zz_stage1Out_payload_wayValid = valid_0_2;
      5'b00011 : _zz_stage1Out_payload_wayValid = valid_0_3;
      5'b00100 : _zz_stage1Out_payload_wayValid = valid_0_4;
      5'b00101 : _zz_stage1Out_payload_wayValid = valid_0_5;
      5'b00110 : _zz_stage1Out_payload_wayValid = valid_0_6;
      5'b00111 : _zz_stage1Out_payload_wayValid = valid_0_7;
      5'b01000 : _zz_stage1Out_payload_wayValid = valid_0_8;
      5'b01001 : _zz_stage1Out_payload_wayValid = valid_0_9;
      5'b01010 : _zz_stage1Out_payload_wayValid = valid_0_10;
      5'b01011 : _zz_stage1Out_payload_wayValid = valid_0_11;
      5'b01100 : _zz_stage1Out_payload_wayValid = valid_0_12;
      5'b01101 : _zz_stage1Out_payload_wayValid = valid_0_13;
      5'b01110 : _zz_stage1Out_payload_wayValid = valid_0_14;
      5'b01111 : _zz_stage1Out_payload_wayValid = valid_0_15;
      5'b10000 : _zz_stage1Out_payload_wayValid = valid_0_16;
      5'b10001 : _zz_stage1Out_payload_wayValid = valid_0_17;
      5'b10010 : _zz_stage1Out_payload_wayValid = valid_0_18;
      5'b10011 : _zz_stage1Out_payload_wayValid = valid_0_19;
      5'b10100 : _zz_stage1Out_payload_wayValid = valid_0_20;
      5'b10101 : _zz_stage1Out_payload_wayValid = valid_0_21;
      5'b10110 : _zz_stage1Out_payload_wayValid = valid_0_22;
      5'b10111 : _zz_stage1Out_payload_wayValid = valid_0_23;
      5'b11000 : _zz_stage1Out_payload_wayValid = valid_0_24;
      5'b11001 : _zz_stage1Out_payload_wayValid = valid_0_25;
      5'b11010 : _zz_stage1Out_payload_wayValid = valid_0_26;
      5'b11011 : _zz_stage1Out_payload_wayValid = valid_0_27;
      5'b11100 : _zz_stage1Out_payload_wayValid = valid_0_28;
      5'b11101 : _zz_stage1Out_payload_wayValid = valid_0_29;
      5'b11110 : _zz_stage1Out_payload_wayValid = valid_0_30;
      default : _zz_stage1Out_payload_wayValid = valid_0_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayDirty_1)
      5'b00000 : _zz_stage1Out_payload_wayDirty = dirty_0_0;
      5'b00001 : _zz_stage1Out_payload_wayDirty = dirty_0_1;
      5'b00010 : _zz_stage1Out_payload_wayDirty = dirty_0_2;
      5'b00011 : _zz_stage1Out_payload_wayDirty = dirty_0_3;
      5'b00100 : _zz_stage1Out_payload_wayDirty = dirty_0_4;
      5'b00101 : _zz_stage1Out_payload_wayDirty = dirty_0_5;
      5'b00110 : _zz_stage1Out_payload_wayDirty = dirty_0_6;
      5'b00111 : _zz_stage1Out_payload_wayDirty = dirty_0_7;
      5'b01000 : _zz_stage1Out_payload_wayDirty = dirty_0_8;
      5'b01001 : _zz_stage1Out_payload_wayDirty = dirty_0_9;
      5'b01010 : _zz_stage1Out_payload_wayDirty = dirty_0_10;
      5'b01011 : _zz_stage1Out_payload_wayDirty = dirty_0_11;
      5'b01100 : _zz_stage1Out_payload_wayDirty = dirty_0_12;
      5'b01101 : _zz_stage1Out_payload_wayDirty = dirty_0_13;
      5'b01110 : _zz_stage1Out_payload_wayDirty = dirty_0_14;
      5'b01111 : _zz_stage1Out_payload_wayDirty = dirty_0_15;
      5'b10000 : _zz_stage1Out_payload_wayDirty = dirty_0_16;
      5'b10001 : _zz_stage1Out_payload_wayDirty = dirty_0_17;
      5'b10010 : _zz_stage1Out_payload_wayDirty = dirty_0_18;
      5'b10011 : _zz_stage1Out_payload_wayDirty = dirty_0_19;
      5'b10100 : _zz_stage1Out_payload_wayDirty = dirty_0_20;
      5'b10101 : _zz_stage1Out_payload_wayDirty = dirty_0_21;
      5'b10110 : _zz_stage1Out_payload_wayDirty = dirty_0_22;
      5'b10111 : _zz_stage1Out_payload_wayDirty = dirty_0_23;
      5'b11000 : _zz_stage1Out_payload_wayDirty = dirty_0_24;
      5'b11001 : _zz_stage1Out_payload_wayDirty = dirty_0_25;
      5'b11010 : _zz_stage1Out_payload_wayDirty = dirty_0_26;
      5'b11011 : _zz_stage1Out_payload_wayDirty = dirty_0_27;
      5'b11100 : _zz_stage1Out_payload_wayDirty = dirty_0_28;
      5'b11101 : _zz_stage1Out_payload_wayDirty = dirty_0_29;
      5'b11110 : _zz_stage1Out_payload_wayDirty = dirty_0_30;
      default : _zz_stage1Out_payload_wayDirty = dirty_0_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_4)
      5'b00000 : _zz_stage1Out_payload_wayValid_3 = valid_1_0;
      5'b00001 : _zz_stage1Out_payload_wayValid_3 = valid_1_1;
      5'b00010 : _zz_stage1Out_payload_wayValid_3 = valid_1_2;
      5'b00011 : _zz_stage1Out_payload_wayValid_3 = valid_1_3;
      5'b00100 : _zz_stage1Out_payload_wayValid_3 = valid_1_4;
      5'b00101 : _zz_stage1Out_payload_wayValid_3 = valid_1_5;
      5'b00110 : _zz_stage1Out_payload_wayValid_3 = valid_1_6;
      5'b00111 : _zz_stage1Out_payload_wayValid_3 = valid_1_7;
      5'b01000 : _zz_stage1Out_payload_wayValid_3 = valid_1_8;
      5'b01001 : _zz_stage1Out_payload_wayValid_3 = valid_1_9;
      5'b01010 : _zz_stage1Out_payload_wayValid_3 = valid_1_10;
      5'b01011 : _zz_stage1Out_payload_wayValid_3 = valid_1_11;
      5'b01100 : _zz_stage1Out_payload_wayValid_3 = valid_1_12;
      5'b01101 : _zz_stage1Out_payload_wayValid_3 = valid_1_13;
      5'b01110 : _zz_stage1Out_payload_wayValid_3 = valid_1_14;
      5'b01111 : _zz_stage1Out_payload_wayValid_3 = valid_1_15;
      5'b10000 : _zz_stage1Out_payload_wayValid_3 = valid_1_16;
      5'b10001 : _zz_stage1Out_payload_wayValid_3 = valid_1_17;
      5'b10010 : _zz_stage1Out_payload_wayValid_3 = valid_1_18;
      5'b10011 : _zz_stage1Out_payload_wayValid_3 = valid_1_19;
      5'b10100 : _zz_stage1Out_payload_wayValid_3 = valid_1_20;
      5'b10101 : _zz_stage1Out_payload_wayValid_3 = valid_1_21;
      5'b10110 : _zz_stage1Out_payload_wayValid_3 = valid_1_22;
      5'b10111 : _zz_stage1Out_payload_wayValid_3 = valid_1_23;
      5'b11000 : _zz_stage1Out_payload_wayValid_3 = valid_1_24;
      5'b11001 : _zz_stage1Out_payload_wayValid_3 = valid_1_25;
      5'b11010 : _zz_stage1Out_payload_wayValid_3 = valid_1_26;
      5'b11011 : _zz_stage1Out_payload_wayValid_3 = valid_1_27;
      5'b11100 : _zz_stage1Out_payload_wayValid_3 = valid_1_28;
      5'b11101 : _zz_stage1Out_payload_wayValid_3 = valid_1_29;
      5'b11110 : _zz_stage1Out_payload_wayValid_3 = valid_1_30;
      default : _zz_stage1Out_payload_wayValid_3 = valid_1_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayDirty_4)
      5'b00000 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_0;
      5'b00001 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_1;
      5'b00010 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_2;
      5'b00011 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_3;
      5'b00100 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_4;
      5'b00101 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_5;
      5'b00110 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_6;
      5'b00111 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_7;
      5'b01000 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_8;
      5'b01001 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_9;
      5'b01010 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_10;
      5'b01011 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_11;
      5'b01100 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_12;
      5'b01101 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_13;
      5'b01110 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_14;
      5'b01111 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_15;
      5'b10000 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_16;
      5'b10001 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_17;
      5'b10010 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_18;
      5'b10011 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_19;
      5'b10100 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_20;
      5'b10101 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_21;
      5'b10110 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_22;
      5'b10111 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_23;
      5'b11000 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_24;
      5'b11001 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_25;
      5'b11010 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_26;
      5'b11011 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_27;
      5'b11100 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_28;
      5'b11101 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_29;
      5'b11110 : _zz_stage1Out_payload_wayDirty_3 = dirty_1_30;
      default : _zz_stage1Out_payload_wayDirty_3 = dirty_1_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_7)
      5'b00000 : _zz_stage1Out_payload_wayValid_6 = valid_2_0;
      5'b00001 : _zz_stage1Out_payload_wayValid_6 = valid_2_1;
      5'b00010 : _zz_stage1Out_payload_wayValid_6 = valid_2_2;
      5'b00011 : _zz_stage1Out_payload_wayValid_6 = valid_2_3;
      5'b00100 : _zz_stage1Out_payload_wayValid_6 = valid_2_4;
      5'b00101 : _zz_stage1Out_payload_wayValid_6 = valid_2_5;
      5'b00110 : _zz_stage1Out_payload_wayValid_6 = valid_2_6;
      5'b00111 : _zz_stage1Out_payload_wayValid_6 = valid_2_7;
      5'b01000 : _zz_stage1Out_payload_wayValid_6 = valid_2_8;
      5'b01001 : _zz_stage1Out_payload_wayValid_6 = valid_2_9;
      5'b01010 : _zz_stage1Out_payload_wayValid_6 = valid_2_10;
      5'b01011 : _zz_stage1Out_payload_wayValid_6 = valid_2_11;
      5'b01100 : _zz_stage1Out_payload_wayValid_6 = valid_2_12;
      5'b01101 : _zz_stage1Out_payload_wayValid_6 = valid_2_13;
      5'b01110 : _zz_stage1Out_payload_wayValid_6 = valid_2_14;
      5'b01111 : _zz_stage1Out_payload_wayValid_6 = valid_2_15;
      5'b10000 : _zz_stage1Out_payload_wayValid_6 = valid_2_16;
      5'b10001 : _zz_stage1Out_payload_wayValid_6 = valid_2_17;
      5'b10010 : _zz_stage1Out_payload_wayValid_6 = valid_2_18;
      5'b10011 : _zz_stage1Out_payload_wayValid_6 = valid_2_19;
      5'b10100 : _zz_stage1Out_payload_wayValid_6 = valid_2_20;
      5'b10101 : _zz_stage1Out_payload_wayValid_6 = valid_2_21;
      5'b10110 : _zz_stage1Out_payload_wayValid_6 = valid_2_22;
      5'b10111 : _zz_stage1Out_payload_wayValid_6 = valid_2_23;
      5'b11000 : _zz_stage1Out_payload_wayValid_6 = valid_2_24;
      5'b11001 : _zz_stage1Out_payload_wayValid_6 = valid_2_25;
      5'b11010 : _zz_stage1Out_payload_wayValid_6 = valid_2_26;
      5'b11011 : _zz_stage1Out_payload_wayValid_6 = valid_2_27;
      5'b11100 : _zz_stage1Out_payload_wayValid_6 = valid_2_28;
      5'b11101 : _zz_stage1Out_payload_wayValid_6 = valid_2_29;
      5'b11110 : _zz_stage1Out_payload_wayValid_6 = valid_2_30;
      default : _zz_stage1Out_payload_wayValid_6 = valid_2_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayDirty_7)
      5'b00000 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_0;
      5'b00001 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_1;
      5'b00010 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_2;
      5'b00011 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_3;
      5'b00100 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_4;
      5'b00101 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_5;
      5'b00110 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_6;
      5'b00111 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_7;
      5'b01000 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_8;
      5'b01001 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_9;
      5'b01010 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_10;
      5'b01011 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_11;
      5'b01100 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_12;
      5'b01101 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_13;
      5'b01110 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_14;
      5'b01111 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_15;
      5'b10000 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_16;
      5'b10001 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_17;
      5'b10010 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_18;
      5'b10011 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_19;
      5'b10100 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_20;
      5'b10101 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_21;
      5'b10110 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_22;
      5'b10111 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_23;
      5'b11000 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_24;
      5'b11001 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_25;
      5'b11010 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_26;
      5'b11011 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_27;
      5'b11100 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_28;
      5'b11101 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_29;
      5'b11110 : _zz_stage1Out_payload_wayDirty_6 = dirty_2_30;
      default : _zz_stage1Out_payload_wayDirty_6 = dirty_2_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_10)
      5'b00000 : _zz_stage1Out_payload_wayValid_9 = valid_3_0;
      5'b00001 : _zz_stage1Out_payload_wayValid_9 = valid_3_1;
      5'b00010 : _zz_stage1Out_payload_wayValid_9 = valid_3_2;
      5'b00011 : _zz_stage1Out_payload_wayValid_9 = valid_3_3;
      5'b00100 : _zz_stage1Out_payload_wayValid_9 = valid_3_4;
      5'b00101 : _zz_stage1Out_payload_wayValid_9 = valid_3_5;
      5'b00110 : _zz_stage1Out_payload_wayValid_9 = valid_3_6;
      5'b00111 : _zz_stage1Out_payload_wayValid_9 = valid_3_7;
      5'b01000 : _zz_stage1Out_payload_wayValid_9 = valid_3_8;
      5'b01001 : _zz_stage1Out_payload_wayValid_9 = valid_3_9;
      5'b01010 : _zz_stage1Out_payload_wayValid_9 = valid_3_10;
      5'b01011 : _zz_stage1Out_payload_wayValid_9 = valid_3_11;
      5'b01100 : _zz_stage1Out_payload_wayValid_9 = valid_3_12;
      5'b01101 : _zz_stage1Out_payload_wayValid_9 = valid_3_13;
      5'b01110 : _zz_stage1Out_payload_wayValid_9 = valid_3_14;
      5'b01111 : _zz_stage1Out_payload_wayValid_9 = valid_3_15;
      5'b10000 : _zz_stage1Out_payload_wayValid_9 = valid_3_16;
      5'b10001 : _zz_stage1Out_payload_wayValid_9 = valid_3_17;
      5'b10010 : _zz_stage1Out_payload_wayValid_9 = valid_3_18;
      5'b10011 : _zz_stage1Out_payload_wayValid_9 = valid_3_19;
      5'b10100 : _zz_stage1Out_payload_wayValid_9 = valid_3_20;
      5'b10101 : _zz_stage1Out_payload_wayValid_9 = valid_3_21;
      5'b10110 : _zz_stage1Out_payload_wayValid_9 = valid_3_22;
      5'b10111 : _zz_stage1Out_payload_wayValid_9 = valid_3_23;
      5'b11000 : _zz_stage1Out_payload_wayValid_9 = valid_3_24;
      5'b11001 : _zz_stage1Out_payload_wayValid_9 = valid_3_25;
      5'b11010 : _zz_stage1Out_payload_wayValid_9 = valid_3_26;
      5'b11011 : _zz_stage1Out_payload_wayValid_9 = valid_3_27;
      5'b11100 : _zz_stage1Out_payload_wayValid_9 = valid_3_28;
      5'b11101 : _zz_stage1Out_payload_wayValid_9 = valid_3_29;
      5'b11110 : _zz_stage1Out_payload_wayValid_9 = valid_3_30;
      default : _zz_stage1Out_payload_wayValid_9 = valid_3_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayDirty_10)
      5'b00000 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_0;
      5'b00001 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_1;
      5'b00010 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_2;
      5'b00011 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_3;
      5'b00100 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_4;
      5'b00101 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_5;
      5'b00110 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_6;
      5'b00111 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_7;
      5'b01000 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_8;
      5'b01001 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_9;
      5'b01010 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_10;
      5'b01011 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_11;
      5'b01100 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_12;
      5'b01101 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_13;
      5'b01110 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_14;
      5'b01111 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_15;
      5'b10000 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_16;
      5'b10001 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_17;
      5'b10010 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_18;
      5'b10011 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_19;
      5'b10100 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_20;
      5'b10101 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_21;
      5'b10110 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_22;
      5'b10111 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_23;
      5'b11000 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_24;
      5'b11001 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_25;
      5'b11010 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_26;
      5'b11011 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_27;
      5'b11100 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_28;
      5'b11101 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_29;
      5'b11110 : _zz_stage1Out_payload_wayDirty_9 = dirty_3_30;
      default : _zz_stage1Out_payload_wayDirty_9 = dirty_3_31;
    endcase
  end

  always @(*) begin
    case(_zz_writeBufferHeadNext_12)
      3'b000 : _zz_writeBufferHeadNext_11 = _zz_writeBufferHeadNext;
      3'b001 : _zz_writeBufferHeadNext_11 = _zz_writeBufferHeadNext_1;
      3'b010 : _zz_writeBufferHeadNext_11 = _zz_writeBufferHeadNext_2;
      3'b011 : _zz_writeBufferHeadNext_11 = _zz_writeBufferHeadNext_3;
      3'b100 : _zz_writeBufferHeadNext_11 = _zz_writeBufferHeadNext_4;
      3'b101 : _zz_writeBufferHeadNext_11 = _zz_writeBufferHeadNext_5;
      3'b110 : _zz_writeBufferHeadNext_11 = _zz_writeBufferHeadNext_6;
      default : _zz_writeBufferHeadNext_11 = _zz_writeBufferHeadNext_7;
    endcase
  end

  always @(*) begin
    case(_zz_writeBufferHeadNext_14)
      3'b000 : _zz_writeBufferHeadNext_13 = _zz_writeBufferHeadNext;
      3'b001 : _zz_writeBufferHeadNext_13 = _zz_writeBufferHeadNext_1;
      3'b010 : _zz_writeBufferHeadNext_13 = _zz_writeBufferHeadNext_2;
      3'b011 : _zz_writeBufferHeadNext_13 = _zz_writeBufferHeadNext_3;
      3'b100 : _zz_writeBufferHeadNext_13 = _zz_writeBufferHeadNext_4;
      3'b101 : _zz_writeBufferHeadNext_13 = _zz_writeBufferHeadNext_5;
      3'b110 : _zz_writeBufferHeadNext_13 = _zz_writeBufferHeadNext_6;
      default : _zz_writeBufferHeadNext_13 = _zz_writeBufferHeadNext_7;
    endcase
  end

  always @(*) begin
    case(_zz_writeBufferHeadNext_16)
      3'b000 : _zz_writeBufferHeadNext_15 = _zz_writeBufferHeadNext;
      3'b001 : _zz_writeBufferHeadNext_15 = _zz_writeBufferHeadNext_1;
      3'b010 : _zz_writeBufferHeadNext_15 = _zz_writeBufferHeadNext_2;
      3'b011 : _zz_writeBufferHeadNext_15 = _zz_writeBufferHeadNext_3;
      3'b100 : _zz_writeBufferHeadNext_15 = _zz_writeBufferHeadNext_4;
      3'b101 : _zz_writeBufferHeadNext_15 = _zz_writeBufferHeadNext_5;
      3'b110 : _zz_writeBufferHeadNext_15 = _zz_writeBufferHeadNext_6;
      default : _zz_writeBufferHeadNext_15 = _zz_writeBufferHeadNext_7;
    endcase
  end

  always @(*) begin
    case(writeBufferTail)
      3'b000 : begin
        _zz__zz_writeBufferAvail = writeBuffer_0_valid;
        _zz_latestWrite_robIdx = writeBuffer_0_robIdx;
        _zz_latestWrite_waySelect = writeBuffer_0_waySelect;
        _zz_latestWrite_prevData = writeBuffer_0_prevData;
        _zz_latestWrite_prevDirty = writeBuffer_0_prevDirty;
        _zz_latestWrite_index = writeBuffer_0_index;
        _zz_latestWrite_miss = writeBuffer_0_miss;
      end
      3'b001 : begin
        _zz__zz_writeBufferAvail = writeBuffer_1_valid;
        _zz_latestWrite_robIdx = writeBuffer_1_robIdx;
        _zz_latestWrite_waySelect = writeBuffer_1_waySelect;
        _zz_latestWrite_prevData = writeBuffer_1_prevData;
        _zz_latestWrite_prevDirty = writeBuffer_1_prevDirty;
        _zz_latestWrite_index = writeBuffer_1_index;
        _zz_latestWrite_miss = writeBuffer_1_miss;
      end
      3'b010 : begin
        _zz__zz_writeBufferAvail = writeBuffer_2_valid;
        _zz_latestWrite_robIdx = writeBuffer_2_robIdx;
        _zz_latestWrite_waySelect = writeBuffer_2_waySelect;
        _zz_latestWrite_prevData = writeBuffer_2_prevData;
        _zz_latestWrite_prevDirty = writeBuffer_2_prevDirty;
        _zz_latestWrite_index = writeBuffer_2_index;
        _zz_latestWrite_miss = writeBuffer_2_miss;
      end
      3'b011 : begin
        _zz__zz_writeBufferAvail = writeBuffer_3_valid;
        _zz_latestWrite_robIdx = writeBuffer_3_robIdx;
        _zz_latestWrite_waySelect = writeBuffer_3_waySelect;
        _zz_latestWrite_prevData = writeBuffer_3_prevData;
        _zz_latestWrite_prevDirty = writeBuffer_3_prevDirty;
        _zz_latestWrite_index = writeBuffer_3_index;
        _zz_latestWrite_miss = writeBuffer_3_miss;
      end
      3'b100 : begin
        _zz__zz_writeBufferAvail = writeBuffer_4_valid;
        _zz_latestWrite_robIdx = writeBuffer_4_robIdx;
        _zz_latestWrite_waySelect = writeBuffer_4_waySelect;
        _zz_latestWrite_prevData = writeBuffer_4_prevData;
        _zz_latestWrite_prevDirty = writeBuffer_4_prevDirty;
        _zz_latestWrite_index = writeBuffer_4_index;
        _zz_latestWrite_miss = writeBuffer_4_miss;
      end
      3'b101 : begin
        _zz__zz_writeBufferAvail = writeBuffer_5_valid;
        _zz_latestWrite_robIdx = writeBuffer_5_robIdx;
        _zz_latestWrite_waySelect = writeBuffer_5_waySelect;
        _zz_latestWrite_prevData = writeBuffer_5_prevData;
        _zz_latestWrite_prevDirty = writeBuffer_5_prevDirty;
        _zz_latestWrite_index = writeBuffer_5_index;
        _zz_latestWrite_miss = writeBuffer_5_miss;
      end
      3'b110 : begin
        _zz__zz_writeBufferAvail = writeBuffer_6_valid;
        _zz_latestWrite_robIdx = writeBuffer_6_robIdx;
        _zz_latestWrite_waySelect = writeBuffer_6_waySelect;
        _zz_latestWrite_prevData = writeBuffer_6_prevData;
        _zz_latestWrite_prevDirty = writeBuffer_6_prevDirty;
        _zz_latestWrite_index = writeBuffer_6_index;
        _zz_latestWrite_miss = writeBuffer_6_miss;
      end
      default : begin
        _zz__zz_writeBufferAvail = writeBuffer_7_valid;
        _zz_latestWrite_robIdx = writeBuffer_7_robIdx;
        _zz_latestWrite_waySelect = writeBuffer_7_waySelect;
        _zz_latestWrite_prevData = writeBuffer_7_prevData;
        _zz_latestWrite_prevDirty = writeBuffer_7_prevDirty;
        _zz_latestWrite_index = writeBuffer_7_index;
        _zz_latestWrite_miss = writeBuffer_7_miss;
      end
    endcase
  end

  always @(*) begin
    case(_zz_io_output_payload_data_2)
      2'b00 : begin
        _zz__zz_writeBuffer_0_prevData = dataRead_0;
        _zz__zz_writeBuffer_0_prevDirty = _zz_missBuffer_0_writeBack;
        _zz_io_output_payload_data_3 = dataShuffle_0;
      end
      2'b01 : begin
        _zz__zz_writeBuffer_0_prevData = dataRead_1;
        _zz__zz_writeBuffer_0_prevDirty = _zz_missBuffer_0_writeBack_1;
        _zz_io_output_payload_data_3 = dataShuffle_1;
      end
      2'b10 : begin
        _zz__zz_writeBuffer_0_prevData = dataRead_2;
        _zz__zz_writeBuffer_0_prevDirty = _zz_missBuffer_0_writeBack_2;
        _zz_io_output_payload_data_3 = dataShuffle_2;
      end
      default : begin
        _zz__zz_writeBuffer_0_prevData = dataRead_3;
        _zz__zz_writeBuffer_0_prevDirty = _zz_missBuffer_0_writeBack_3;
        _zz_io_output_payload_data_3 = dataShuffle_3;
      end
    endcase
  end

  always @(*) begin
    case(_zz_missBuffer_0_writeBack_7)
      2'b00 : begin
        _zz_missBuffer_0_writeBack_8 = _zz_missBuffer_0_writeBack;
        _zz_missBuffer_0_prevPaddr = tagRead_0;
      end
      2'b01 : begin
        _zz_missBuffer_0_writeBack_8 = _zz_missBuffer_0_writeBack_1;
        _zz_missBuffer_0_prevPaddr = tagRead_1;
      end
      2'b10 : begin
        _zz_missBuffer_0_writeBack_8 = _zz_missBuffer_0_writeBack_2;
        _zz_missBuffer_0_prevPaddr = tagRead_2;
      end
      default : begin
        _zz_missBuffer_0_writeBack_8 = _zz_missBuffer_0_writeBack_3;
        _zz_missBuffer_0_prevPaddr = tagRead_3;
      end
    endcase
  end

  always @(*) begin
    case(_zz_io_axi_wdata_3)
      2'b00 : _zz_io_axi_wdata_2 = portRData1_0;
      2'b01 : _zz_io_axi_wdata_2 = portRData1_1;
      2'b10 : _zz_io_axi_wdata_2 = portRData1_2;
      default : _zz_io_axi_wdata_2 = portRData1_3;
    endcase
  end

  always @(*) begin
    case(_zz_cacopPAddr_1)
      2'b00 : _zz_cacopPAddr = tagRead_0;
      2'b01 : _zz_cacopPAddr = tagRead_1;
      2'b10 : _zz_cacopPAddr = tagRead_2;
      default : _zz_cacopPAddr = tagRead_3;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_1)
      5'b00000 : _zz__zz_wayToReplace = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace = lruBit_30_0;
      default : _zz__zz_wayToReplace = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_3)
      5'b00000 : _zz__zz_wayToReplace_2 = lruBit_0_1;
      5'b00001 : _zz__zz_wayToReplace_2 = lruBit_1_1;
      5'b00010 : _zz__zz_wayToReplace_2 = lruBit_2_1;
      5'b00011 : _zz__zz_wayToReplace_2 = lruBit_3_1;
      5'b00100 : _zz__zz_wayToReplace_2 = lruBit_4_1;
      5'b00101 : _zz__zz_wayToReplace_2 = lruBit_5_1;
      5'b00110 : _zz__zz_wayToReplace_2 = lruBit_6_1;
      5'b00111 : _zz__zz_wayToReplace_2 = lruBit_7_1;
      5'b01000 : _zz__zz_wayToReplace_2 = lruBit_8_1;
      5'b01001 : _zz__zz_wayToReplace_2 = lruBit_9_1;
      5'b01010 : _zz__zz_wayToReplace_2 = lruBit_10_1;
      5'b01011 : _zz__zz_wayToReplace_2 = lruBit_11_1;
      5'b01100 : _zz__zz_wayToReplace_2 = lruBit_12_1;
      5'b01101 : _zz__zz_wayToReplace_2 = lruBit_13_1;
      5'b01110 : _zz__zz_wayToReplace_2 = lruBit_14_1;
      5'b01111 : _zz__zz_wayToReplace_2 = lruBit_15_1;
      5'b10000 : _zz__zz_wayToReplace_2 = lruBit_16_1;
      5'b10001 : _zz__zz_wayToReplace_2 = lruBit_17_1;
      5'b10010 : _zz__zz_wayToReplace_2 = lruBit_18_1;
      5'b10011 : _zz__zz_wayToReplace_2 = lruBit_19_1;
      5'b10100 : _zz__zz_wayToReplace_2 = lruBit_20_1;
      5'b10101 : _zz__zz_wayToReplace_2 = lruBit_21_1;
      5'b10110 : _zz__zz_wayToReplace_2 = lruBit_22_1;
      5'b10111 : _zz__zz_wayToReplace_2 = lruBit_23_1;
      5'b11000 : _zz__zz_wayToReplace_2 = lruBit_24_1;
      5'b11001 : _zz__zz_wayToReplace_2 = lruBit_25_1;
      5'b11010 : _zz__zz_wayToReplace_2 = lruBit_26_1;
      5'b11011 : _zz__zz_wayToReplace_2 = lruBit_27_1;
      5'b11100 : _zz__zz_wayToReplace_2 = lruBit_28_1;
      5'b11101 : _zz__zz_wayToReplace_2 = lruBit_29_1;
      5'b11110 : _zz__zz_wayToReplace_2 = lruBit_30_1;
      default : _zz__zz_wayToReplace_2 = lruBit_31_1;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_1_2)
      5'b00000 : _zz__zz_wayToReplace_1_1 = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace_1_1 = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace_1_1 = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace_1_1 = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace_1_1 = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace_1_1 = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace_1_1 = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace_1_1 = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace_1_1 = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace_1_1 = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace_1_1 = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace_1_1 = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace_1_1 = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace_1_1 = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace_1_1 = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace_1_1 = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace_1_1 = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace_1_1 = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace_1_1 = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace_1_1 = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace_1_1 = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace_1_1 = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace_1_1 = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace_1_1 = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace_1_1 = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace_1_1 = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace_1_1 = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace_1_1 = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace_1_1 = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace_1_1 = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace_1_1 = lruBit_30_0;
      default : _zz__zz_wayToReplace_1_1 = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_1_4)
      5'b00000 : _zz__zz_wayToReplace_1_3 = lruBit_0_1;
      5'b00001 : _zz__zz_wayToReplace_1_3 = lruBit_1_1;
      5'b00010 : _zz__zz_wayToReplace_1_3 = lruBit_2_1;
      5'b00011 : _zz__zz_wayToReplace_1_3 = lruBit_3_1;
      5'b00100 : _zz__zz_wayToReplace_1_3 = lruBit_4_1;
      5'b00101 : _zz__zz_wayToReplace_1_3 = lruBit_5_1;
      5'b00110 : _zz__zz_wayToReplace_1_3 = lruBit_6_1;
      5'b00111 : _zz__zz_wayToReplace_1_3 = lruBit_7_1;
      5'b01000 : _zz__zz_wayToReplace_1_3 = lruBit_8_1;
      5'b01001 : _zz__zz_wayToReplace_1_3 = lruBit_9_1;
      5'b01010 : _zz__zz_wayToReplace_1_3 = lruBit_10_1;
      5'b01011 : _zz__zz_wayToReplace_1_3 = lruBit_11_1;
      5'b01100 : _zz__zz_wayToReplace_1_3 = lruBit_12_1;
      5'b01101 : _zz__zz_wayToReplace_1_3 = lruBit_13_1;
      5'b01110 : _zz__zz_wayToReplace_1_3 = lruBit_14_1;
      5'b01111 : _zz__zz_wayToReplace_1_3 = lruBit_15_1;
      5'b10000 : _zz__zz_wayToReplace_1_3 = lruBit_16_1;
      5'b10001 : _zz__zz_wayToReplace_1_3 = lruBit_17_1;
      5'b10010 : _zz__zz_wayToReplace_1_3 = lruBit_18_1;
      5'b10011 : _zz__zz_wayToReplace_1_3 = lruBit_19_1;
      5'b10100 : _zz__zz_wayToReplace_1_3 = lruBit_20_1;
      5'b10101 : _zz__zz_wayToReplace_1_3 = lruBit_21_1;
      5'b10110 : _zz__zz_wayToReplace_1_3 = lruBit_22_1;
      5'b10111 : _zz__zz_wayToReplace_1_3 = lruBit_23_1;
      5'b11000 : _zz__zz_wayToReplace_1_3 = lruBit_24_1;
      5'b11001 : _zz__zz_wayToReplace_1_3 = lruBit_25_1;
      5'b11010 : _zz__zz_wayToReplace_1_3 = lruBit_26_1;
      5'b11011 : _zz__zz_wayToReplace_1_3 = lruBit_27_1;
      5'b11100 : _zz__zz_wayToReplace_1_3 = lruBit_28_1;
      5'b11101 : _zz__zz_wayToReplace_1_3 = lruBit_29_1;
      5'b11110 : _zz__zz_wayToReplace_1_3 = lruBit_30_1;
      default : _zz__zz_wayToReplace_1_3 = lruBit_31_1;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_2_2)
      5'b00000 : _zz__zz_wayToReplace_2_1 = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace_2_1 = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace_2_1 = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace_2_1 = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace_2_1 = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace_2_1 = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace_2_1 = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace_2_1 = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace_2_1 = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace_2_1 = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace_2_1 = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace_2_1 = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace_2_1 = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace_2_1 = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace_2_1 = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace_2_1 = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace_2_1 = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace_2_1 = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace_2_1 = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace_2_1 = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace_2_1 = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace_2_1 = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace_2_1 = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace_2_1 = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace_2_1 = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace_2_1 = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace_2_1 = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace_2_1 = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace_2_1 = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace_2_1 = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace_2_1 = lruBit_30_0;
      default : _zz__zz_wayToReplace_2_1 = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_2_4)
      5'b00000 : _zz__zz_wayToReplace_2_3 = lruBit_0_2;
      5'b00001 : _zz__zz_wayToReplace_2_3 = lruBit_1_2;
      5'b00010 : _zz__zz_wayToReplace_2_3 = lruBit_2_2;
      5'b00011 : _zz__zz_wayToReplace_2_3 = lruBit_3_2;
      5'b00100 : _zz__zz_wayToReplace_2_3 = lruBit_4_2;
      5'b00101 : _zz__zz_wayToReplace_2_3 = lruBit_5_2;
      5'b00110 : _zz__zz_wayToReplace_2_3 = lruBit_6_2;
      5'b00111 : _zz__zz_wayToReplace_2_3 = lruBit_7_2;
      5'b01000 : _zz__zz_wayToReplace_2_3 = lruBit_8_2;
      5'b01001 : _zz__zz_wayToReplace_2_3 = lruBit_9_2;
      5'b01010 : _zz__zz_wayToReplace_2_3 = lruBit_10_2;
      5'b01011 : _zz__zz_wayToReplace_2_3 = lruBit_11_2;
      5'b01100 : _zz__zz_wayToReplace_2_3 = lruBit_12_2;
      5'b01101 : _zz__zz_wayToReplace_2_3 = lruBit_13_2;
      5'b01110 : _zz__zz_wayToReplace_2_3 = lruBit_14_2;
      5'b01111 : _zz__zz_wayToReplace_2_3 = lruBit_15_2;
      5'b10000 : _zz__zz_wayToReplace_2_3 = lruBit_16_2;
      5'b10001 : _zz__zz_wayToReplace_2_3 = lruBit_17_2;
      5'b10010 : _zz__zz_wayToReplace_2_3 = lruBit_18_2;
      5'b10011 : _zz__zz_wayToReplace_2_3 = lruBit_19_2;
      5'b10100 : _zz__zz_wayToReplace_2_3 = lruBit_20_2;
      5'b10101 : _zz__zz_wayToReplace_2_3 = lruBit_21_2;
      5'b10110 : _zz__zz_wayToReplace_2_3 = lruBit_22_2;
      5'b10111 : _zz__zz_wayToReplace_2_3 = lruBit_23_2;
      5'b11000 : _zz__zz_wayToReplace_2_3 = lruBit_24_2;
      5'b11001 : _zz__zz_wayToReplace_2_3 = lruBit_25_2;
      5'b11010 : _zz__zz_wayToReplace_2_3 = lruBit_26_2;
      5'b11011 : _zz__zz_wayToReplace_2_3 = lruBit_27_2;
      5'b11100 : _zz__zz_wayToReplace_2_3 = lruBit_28_2;
      5'b11101 : _zz__zz_wayToReplace_2_3 = lruBit_29_2;
      5'b11110 : _zz__zz_wayToReplace_2_3 = lruBit_30_2;
      default : _zz__zz_wayToReplace_2_3 = lruBit_31_2;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_3_2)
      5'b00000 : _zz__zz_wayToReplace_3_1 = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace_3_1 = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace_3_1 = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace_3_1 = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace_3_1 = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace_3_1 = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace_3_1 = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace_3_1 = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace_3_1 = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace_3_1 = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace_3_1 = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace_3_1 = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace_3_1 = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace_3_1 = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace_3_1 = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace_3_1 = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace_3_1 = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace_3_1 = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace_3_1 = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace_3_1 = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace_3_1 = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace_3_1 = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace_3_1 = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace_3_1 = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace_3_1 = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace_3_1 = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace_3_1 = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace_3_1 = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace_3_1 = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace_3_1 = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace_3_1 = lruBit_30_0;
      default : _zz__zz_wayToReplace_3_1 = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_3_4)
      5'b00000 : _zz__zz_wayToReplace_3_3 = lruBit_0_2;
      5'b00001 : _zz__zz_wayToReplace_3_3 = lruBit_1_2;
      5'b00010 : _zz__zz_wayToReplace_3_3 = lruBit_2_2;
      5'b00011 : _zz__zz_wayToReplace_3_3 = lruBit_3_2;
      5'b00100 : _zz__zz_wayToReplace_3_3 = lruBit_4_2;
      5'b00101 : _zz__zz_wayToReplace_3_3 = lruBit_5_2;
      5'b00110 : _zz__zz_wayToReplace_3_3 = lruBit_6_2;
      5'b00111 : _zz__zz_wayToReplace_3_3 = lruBit_7_2;
      5'b01000 : _zz__zz_wayToReplace_3_3 = lruBit_8_2;
      5'b01001 : _zz__zz_wayToReplace_3_3 = lruBit_9_2;
      5'b01010 : _zz__zz_wayToReplace_3_3 = lruBit_10_2;
      5'b01011 : _zz__zz_wayToReplace_3_3 = lruBit_11_2;
      5'b01100 : _zz__zz_wayToReplace_3_3 = lruBit_12_2;
      5'b01101 : _zz__zz_wayToReplace_3_3 = lruBit_13_2;
      5'b01110 : _zz__zz_wayToReplace_3_3 = lruBit_14_2;
      5'b01111 : _zz__zz_wayToReplace_3_3 = lruBit_15_2;
      5'b10000 : _zz__zz_wayToReplace_3_3 = lruBit_16_2;
      5'b10001 : _zz__zz_wayToReplace_3_3 = lruBit_17_2;
      5'b10010 : _zz__zz_wayToReplace_3_3 = lruBit_18_2;
      5'b10011 : _zz__zz_wayToReplace_3_3 = lruBit_19_2;
      5'b10100 : _zz__zz_wayToReplace_3_3 = lruBit_20_2;
      5'b10101 : _zz__zz_wayToReplace_3_3 = lruBit_21_2;
      5'b10110 : _zz__zz_wayToReplace_3_3 = lruBit_22_2;
      5'b10111 : _zz__zz_wayToReplace_3_3 = lruBit_23_2;
      5'b11000 : _zz__zz_wayToReplace_3_3 = lruBit_24_2;
      5'b11001 : _zz__zz_wayToReplace_3_3 = lruBit_25_2;
      5'b11010 : _zz__zz_wayToReplace_3_3 = lruBit_26_2;
      5'b11011 : _zz__zz_wayToReplace_3_3 = lruBit_27_2;
      5'b11100 : _zz__zz_wayToReplace_3_3 = lruBit_28_2;
      5'b11101 : _zz__zz_wayToReplace_3_3 = lruBit_29_2;
      5'b11110 : _zz__zz_wayToReplace_3_3 = lruBit_30_2;
      default : _zz__zz_wayToReplace_3_3 = lruBit_31_2;
    endcase
  end

  always @(*) begin
    case(writeBufferHeadNext)
      3'b000 : _zz_when_LSU_l567 = writeBuffer_0_valid;
      3'b001 : _zz_when_LSU_l567 = writeBuffer_1_valid;
      3'b010 : _zz_when_LSU_l567 = writeBuffer_2_valid;
      3'b011 : _zz_when_LSU_l567 = writeBuffer_3_valid;
      3'b100 : _zz_when_LSU_l567 = writeBuffer_4_valid;
      3'b101 : _zz_when_LSU_l567 = writeBuffer_5_valid;
      3'b110 : _zz_when_LSU_l567 = writeBuffer_6_valid;
      default : _zz_when_LSU_l567 = writeBuffer_7_valid;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_uop_lsuOp)
      LSUOp_cacop : io_input_payload_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : io_input_payload_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : io_input_payload_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : io_input_payload_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : io_input_payload_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : io_input_payload_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : io_input_payload_uop_lsuOp_string = "ll     ";
      LSUOp_sc : io_input_payload_uop_lsuOp_string = "sc     ";
      LSUOp_ld : io_input_payload_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : io_input_payload_uop_lsuOp_string = "ldu    ";
      LSUOp_st : io_input_payload_uop_lsuOp_string = "st     ";
      LSUOp_preld : io_input_payload_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : io_input_payload_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : io_input_payload_uop_lsuOp_string = "ibar   ";
      default : io_input_payload_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_specialOpBufferUpdate_payload_uop_lsuOp)
      LSUOp_cacop : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "ll     ";
      LSUOp_sc : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "sc     ";
      LSUOp_ld : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "ldu    ";
      LSUOp_st : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "st     ";
      LSUOp_preld : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "ibar   ";
      default : io_specialOpBufferUpdate_payload_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_BOOT : axiCtrl_stateReg_string = "BOOT     ";
      axiCtrl_enumDef_idle : axiCtrl_stateReg_string = "idle     ";
      axiCtrl_enumDef_readReq : axiCtrl_stateReg_string = "readReq  ";
      axiCtrl_enumDef_readFirst : axiCtrl_stateReg_string = "readFirst";
      axiCtrl_enumDef_read : axiCtrl_stateReg_string = "read     ";
      axiCtrl_enumDef_writeReq : axiCtrl_stateReg_string = "writeReq ";
      axiCtrl_enumDef_write : axiCtrl_stateReg_string = "write    ";
      default : axiCtrl_stateReg_string = "?????????";
    endcase
  end
  always @(*) begin
    case(axiCtrl_stateNext)
      axiCtrl_enumDef_BOOT : axiCtrl_stateNext_string = "BOOT     ";
      axiCtrl_enumDef_idle : axiCtrl_stateNext_string = "idle     ";
      axiCtrl_enumDef_readReq : axiCtrl_stateNext_string = "readReq  ";
      axiCtrl_enumDef_readFirst : axiCtrl_stateNext_string = "readFirst";
      axiCtrl_enumDef_read : axiCtrl_stateNext_string = "read     ";
      axiCtrl_enumDef_writeReq : axiCtrl_stateNext_string = "writeReq ";
      axiCtrl_enumDef_write : axiCtrl_stateNext_string = "write    ";
      default : axiCtrl_stateNext_string = "?????????";
    endcase
  end
  always @(*) begin
    case(rollbackCtrl_stateReg)
      rollbackCtrl_enumDef_BOOT : rollbackCtrl_stateReg_string = "BOOT    ";
      rollbackCtrl_enumDef_idle : rollbackCtrl_stateReg_string = "idle    ";
      rollbackCtrl_enumDef_rollback : rollbackCtrl_stateReg_string = "rollback";
      default : rollbackCtrl_stateReg_string = "????????";
    endcase
  end
  always @(*) begin
    case(rollbackCtrl_stateNext)
      rollbackCtrl_enumDef_BOOT : rollbackCtrl_stateNext_string = "BOOT    ";
      rollbackCtrl_enumDef_idle : rollbackCtrl_stateNext_string = "idle    ";
      rollbackCtrl_enumDef_rollback : rollbackCtrl_stateNext_string = "rollback";
      default : rollbackCtrl_stateNext_string = "????????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_wr_en = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
      end
      axiCtrl_enumDef_readReq : begin
        if(when_LSU_l471) begin
          if(when_LSU_l473_3) begin
            _zz_wr_en = 1'b1;
          end
        end
      end
      axiCtrl_enumDef_readFirst : begin
      end
      axiCtrl_enumDef_read : begin
      end
      axiCtrl_enumDef_writeReq : begin
      end
      axiCtrl_enumDef_write : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_wr_en_1 = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
      end
      axiCtrl_enumDef_readReq : begin
        if(when_LSU_l471) begin
          if(when_LSU_l473_2) begin
            _zz_wr_en_1 = 1'b1;
          end
        end
      end
      axiCtrl_enumDef_readFirst : begin
      end
      axiCtrl_enumDef_read : begin
      end
      axiCtrl_enumDef_writeReq : begin
      end
      axiCtrl_enumDef_write : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_wr_en_2 = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
      end
      axiCtrl_enumDef_readReq : begin
        if(when_LSU_l471) begin
          if(when_LSU_l473_1) begin
            _zz_wr_en_2 = 1'b1;
          end
        end
      end
      axiCtrl_enumDef_readFirst : begin
      end
      axiCtrl_enumDef_read : begin
      end
      axiCtrl_enumDef_writeReq : begin
      end
      axiCtrl_enumDef_write : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_wr_en_3 = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
      end
      axiCtrl_enumDef_readReq : begin
        if(when_LSU_l471) begin
          if(when_LSU_l473) begin
            _zz_wr_en_3 = 1'b1;
          end
        end
      end
      axiCtrl_enumDef_readFirst : begin
      end
      axiCtrl_enumDef_read : begin
      end
      axiCtrl_enumDef_writeReq : begin
      end
      axiCtrl_enumDef_write : begin
      end
      default : begin
      end
    endcase
  end

  assign address = (io_input_payload_src1 + io_input_payload_src2);
  assign cacopEn = ((io_ctrl_cacopStoreTag || io_ctrl_cacopIndexInvalidate) || io_ctrl_cacopHitInvalidate);
  always @(*) begin
    stage1Out_thrown_valid = stage1Out_valid;
    if(io_flush) begin
      stage1Out_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    stage1Out_ready = stage1Out_thrown_ready;
    if(io_flush) begin
      stage1Out_ready = 1'b1;
    end
  end

  assign stage1Out_thrown_payload_robIdx = stage1Out_payload_robIdx;
  assign stage1Out_thrown_payload_prd = stage1Out_payload_prd;
  assign stage1Out_thrown_payload_branchResult_targetPC = stage1Out_payload_branchResult_targetPC;
  assign stage1Out_thrown_payload_branchResult_branchResult = stage1Out_payload_branchResult_branchResult;
  assign stage1Out_thrown_payload_branchResult_predictFail = stage1Out_payload_branchResult_predictFail;
  assign stage1Out_thrown_payload_exceptionInfo_exception = stage1Out_payload_exceptionInfo_exception;
  assign stage1Out_thrown_payload_exceptionInfo_eCode = stage1Out_payload_exceptionInfo_eCode;
  assign stage1Out_thrown_payload_exceptionInfo_eSubCode = stage1Out_payload_exceptionInfo_eSubCode;
  assign stage1Out_thrown_payload_storeData = stage1Out_payload_storeData;
  assign stage1Out_thrown_payload_lsCtrlBundle_load = stage1Out_payload_lsCtrlBundle_load;
  assign stage1Out_thrown_payload_lsCtrlBundle_store = stage1Out_payload_lsCtrlBundle_store;
  assign stage1Out_thrown_payload_lsCtrlBundle_signed = stage1Out_payload_lsCtrlBundle_signed;
  assign stage1Out_thrown_payload_lsCtrlBundle_ll = stage1Out_payload_lsCtrlBundle_ll;
  assign stage1Out_thrown_payload_lsCtrlBundle_sc = stage1Out_payload_lsCtrlBundle_sc;
  assign stage1Out_thrown_payload_lsCtrlBundle_lsMask = stage1Out_payload_lsCtrlBundle_lsMask;
  assign stage1Out_thrown_payload_lsCtrlBundle_size = stage1Out_payload_lsCtrlBundle_size;
  assign stage1Out_thrown_payload_lsCtrlBundle_normalMemOp = stage1Out_payload_lsCtrlBundle_normalMemOp;
  assign stage1Out_thrown_payload_vaddr = stage1Out_payload_vaddr;
  assign stage1Out_thrown_payload_tlb_hit = stage1Out_payload_tlb_hit;
  assign stage1Out_thrown_payload_tlb_pageInfo_ppn = stage1Out_payload_tlb_pageInfo_ppn;
  assign stage1Out_thrown_payload_tlb_pageInfo_plv = stage1Out_payload_tlb_pageInfo_plv;
  assign stage1Out_thrown_payload_tlb_pageInfo_mat = stage1Out_payload_tlb_pageInfo_mat;
  assign stage1Out_thrown_payload_tlb_pageInfo_d = stage1Out_payload_tlb_pageInfo_d;
  assign stage1Out_thrown_payload_tlb_pageInfo_v = stage1Out_payload_tlb_pageInfo_v;
  assign stage1Out_thrown_payload_wayValid = stage1Out_payload_wayValid;
  assign stage1Out_thrown_payload_wayDirty = stage1Out_payload_wayDirty;
  assign stage1Out_thrown_payload_isStoreTag = stage1Out_payload_isStoreTag;
  assign stage1Out_thrown_payload_isIndexInvalidate = stage1Out_payload_isIndexInvalidate;
  assign stage1Out_thrown_payload_isHitInvalidate = stage1Out_payload_isHitInvalidate;
  assign stage1Out_thrown_payload_checkTLBException = stage1Out_payload_checkTLBException;
  assign stage1Out_thrown_payload_lsException = stage1Out_payload_lsException;
  always @(*) begin
    stage1Out_thrown_ready = stage1Out_thrown_m2sPipe_ready;
    if(when_Stream_l369) begin
      stage1Out_thrown_ready = 1'b1;
    end
  end

  assign when_Stream_l369 = (! stage1Out_thrown_m2sPipe_valid);
  assign stage1Out_thrown_m2sPipe_valid = stage1Out_thrown_rValid;
  assign stage1Out_thrown_m2sPipe_payload_robIdx = stage1Out_thrown_rData_robIdx;
  assign stage1Out_thrown_m2sPipe_payload_prd = stage1Out_thrown_rData_prd;
  assign stage1Out_thrown_m2sPipe_payload_branchResult_targetPC = stage1Out_thrown_rData_branchResult_targetPC;
  assign stage1Out_thrown_m2sPipe_payload_branchResult_branchResult = stage1Out_thrown_rData_branchResult_branchResult;
  assign stage1Out_thrown_m2sPipe_payload_branchResult_predictFail = stage1Out_thrown_rData_branchResult_predictFail;
  assign stage1Out_thrown_m2sPipe_payload_exceptionInfo_exception = stage1Out_thrown_rData_exceptionInfo_exception;
  assign stage1Out_thrown_m2sPipe_payload_exceptionInfo_eCode = stage1Out_thrown_rData_exceptionInfo_eCode;
  assign stage1Out_thrown_m2sPipe_payload_exceptionInfo_eSubCode = stage1Out_thrown_rData_exceptionInfo_eSubCode;
  assign stage1Out_thrown_m2sPipe_payload_storeData = stage1Out_thrown_rData_storeData;
  assign stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_load = stage1Out_thrown_rData_lsCtrlBundle_load;
  assign stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_store = stage1Out_thrown_rData_lsCtrlBundle_store;
  assign stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_signed = stage1Out_thrown_rData_lsCtrlBundle_signed;
  assign stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_ll = stage1Out_thrown_rData_lsCtrlBundle_ll;
  assign stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_sc = stage1Out_thrown_rData_lsCtrlBundle_sc;
  assign stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_lsMask = stage1Out_thrown_rData_lsCtrlBundle_lsMask;
  assign stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_size = stage1Out_thrown_rData_lsCtrlBundle_size;
  assign stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_normalMemOp = stage1Out_thrown_rData_lsCtrlBundle_normalMemOp;
  assign stage1Out_thrown_m2sPipe_payload_vaddr = stage1Out_thrown_rData_vaddr;
  assign stage1Out_thrown_m2sPipe_payload_tlb_hit = stage1Out_thrown_rData_tlb_hit;
  assign stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_ppn = stage1Out_thrown_rData_tlb_pageInfo_ppn;
  assign stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_plv = stage1Out_thrown_rData_tlb_pageInfo_plv;
  assign stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_mat = stage1Out_thrown_rData_tlb_pageInfo_mat;
  assign stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_d = stage1Out_thrown_rData_tlb_pageInfo_d;
  assign stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_v = stage1Out_thrown_rData_tlb_pageInfo_v;
  assign stage1Out_thrown_m2sPipe_payload_wayValid = stage1Out_thrown_rData_wayValid;
  assign stage1Out_thrown_m2sPipe_payload_wayDirty = stage1Out_thrown_rData_wayDirty;
  assign stage1Out_thrown_m2sPipe_payload_isStoreTag = stage1Out_thrown_rData_isStoreTag;
  assign stage1Out_thrown_m2sPipe_payload_isIndexInvalidate = stage1Out_thrown_rData_isIndexInvalidate;
  assign stage1Out_thrown_m2sPipe_payload_isHitInvalidate = stage1Out_thrown_rData_isHitInvalidate;
  assign stage1Out_thrown_m2sPipe_payload_checkTLBException = stage1Out_thrown_rData_checkTLBException;
  assign stage1Out_thrown_m2sPipe_payload_lsException = stage1Out_thrown_rData_lsException;
  assign stage2In_valid = stage1Out_thrown_m2sPipe_valid;
  assign stage1Out_thrown_m2sPipe_ready = stage2In_ready;
  assign stage2In_payload_robIdx = stage1Out_thrown_m2sPipe_payload_robIdx;
  assign stage2In_payload_prd = stage1Out_thrown_m2sPipe_payload_prd;
  assign stage2In_payload_branchResult_targetPC = stage1Out_thrown_m2sPipe_payload_branchResult_targetPC;
  assign stage2In_payload_branchResult_branchResult = stage1Out_thrown_m2sPipe_payload_branchResult_branchResult;
  assign stage2In_payload_branchResult_predictFail = stage1Out_thrown_m2sPipe_payload_branchResult_predictFail;
  assign stage2In_payload_exceptionInfo_exception = stage1Out_thrown_m2sPipe_payload_exceptionInfo_exception;
  assign stage2In_payload_exceptionInfo_eCode = stage1Out_thrown_m2sPipe_payload_exceptionInfo_eCode;
  assign stage2In_payload_exceptionInfo_eSubCode = stage1Out_thrown_m2sPipe_payload_exceptionInfo_eSubCode;
  assign stage2In_payload_storeData = stage1Out_thrown_m2sPipe_payload_storeData;
  assign stage2In_payload_lsCtrlBundle_load = stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_load;
  assign stage2In_payload_lsCtrlBundle_store = stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_store;
  assign stage2In_payload_lsCtrlBundle_signed = stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_signed;
  assign stage2In_payload_lsCtrlBundle_ll = stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_ll;
  assign stage2In_payload_lsCtrlBundle_sc = stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_sc;
  assign stage2In_payload_lsCtrlBundle_lsMask = stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_lsMask;
  assign stage2In_payload_lsCtrlBundle_size = stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_size;
  assign stage2In_payload_lsCtrlBundle_normalMemOp = stage1Out_thrown_m2sPipe_payload_lsCtrlBundle_normalMemOp;
  assign stage2In_payload_vaddr = stage1Out_thrown_m2sPipe_payload_vaddr;
  assign stage2In_payload_tlb_hit = stage1Out_thrown_m2sPipe_payload_tlb_hit;
  assign stage2In_payload_tlb_pageInfo_ppn = stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_ppn;
  assign stage2In_payload_tlb_pageInfo_plv = stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_plv;
  assign stage2In_payload_tlb_pageInfo_mat = stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_mat;
  assign stage2In_payload_tlb_pageInfo_d = stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_d;
  assign stage2In_payload_tlb_pageInfo_v = stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_v;
  assign stage2In_payload_wayValid = stage1Out_thrown_m2sPipe_payload_wayValid;
  assign stage2In_payload_wayDirty = stage1Out_thrown_m2sPipe_payload_wayDirty;
  assign stage2In_payload_isStoreTag = stage1Out_thrown_m2sPipe_payload_isStoreTag;
  assign stage2In_payload_isIndexInvalidate = stage1Out_thrown_m2sPipe_payload_isIndexInvalidate;
  assign stage2In_payload_isHitInvalidate = stage1Out_thrown_m2sPipe_payload_isHitInvalidate;
  assign stage2In_payload_checkTLBException = stage1Out_thrown_m2sPipe_payload_checkTLBException;
  assign stage2In_payload_lsException = stage1Out_thrown_m2sPipe_payload_lsException;
  assign stage1Out_valid = ((io_input_valid && (! stall)) || cacopEn);
  assign preShiftSize = address[1 : 0];
  assign io_tlb_virtPageNumber = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA[31 : 12] : address[31 : 12]);
  assign io_input_ready = ((stage1Out_ready && (! stall)) || io_flush);
  assign stage1Out_payload_tlb_hit = io_tlb_hit;
  assign stage1Out_payload_tlb_pageInfo_ppn = io_tlb_pageInfo_ppn;
  assign stage1Out_payload_tlb_pageInfo_plv = io_tlb_pageInfo_plv;
  assign stage1Out_payload_tlb_pageInfo_mat = io_tlb_pageInfo_mat;
  assign stage1Out_payload_tlb_pageInfo_d = io_tlb_pageInfo_d;
  assign stage1Out_payload_tlb_pageInfo_v = io_tlb_pageInfo_v;
  assign stage1Out_payload_isStoreTag = io_ctrl_cacopStoreTag;
  assign stage1Out_payload_isIndexInvalidate = io_ctrl_cacopIndexInvalidate;
  assign stage1Out_payload_isHitInvalidate = io_ctrl_cacopHitInvalidate;
  assign stage1Out_payload_robIdx = io_input_payload_robIdx;
  assign stage1Out_payload_prd = io_input_payload_prd;
  assign stage1Out_payload_branchResult_targetPC = io_input_payload_branchResult_targetPC;
  assign stage1Out_payload_branchResult_branchResult = io_input_payload_branchResult_branchResult;
  assign stage1Out_payload_branchResult_predictFail = io_input_payload_branchResult_predictFail;
  assign stage1Out_payload_exceptionInfo_exception = (io_input_payload_exceptionInfo_exception ? io_input_payload_exceptionInfo_exception : exceptionInfo1_exception);
  assign stage1Out_payload_exceptionInfo_eCode = (io_input_payload_exceptionInfo_exception ? io_input_payload_exceptionInfo_eCode : exceptionInfo1_eCode);
  assign stage1Out_payload_exceptionInfo_eSubCode = (io_input_payload_exceptionInfo_exception ? io_input_payload_exceptionInfo_eSubCode : exceptionInfo1_eSubCode);
  assign stage1Out_payload_storeData = _zz_stage1Out_payload_storeData;
  assign stage1Out_payload_vaddr = (cacopEn ? io_ctrl_cacopVA : address);
  assign stage1Out_payload_lsCtrlBundle_load = (((io_input_payload_uop_lsuOp == LSUOp_ld) || (io_input_payload_uop_lsuOp == LSUOp_ldu)) || (io_input_payload_uop_lsuOp == LSUOp_ll));
  assign stage1Out_payload_lsCtrlBundle_store = ((io_input_payload_uop_lsuOp == LSUOp_st) || (io_input_payload_uop_lsuOp == LSUOp_sc));
  assign stage1Out_payload_lsCtrlBundle_signed = (io_input_payload_uop_lsuOp == LSUOp_ld);
  assign stage1Out_payload_lsCtrlBundle_ll = (io_input_payload_uop_lsuOp == LSUOp_ll);
  assign stage1Out_payload_lsCtrlBundle_sc = (io_input_payload_uop_lsuOp == LSUOp_sc);
  assign stage1Out_payload_lsCtrlBundle_lsMask = (io_input_payload_uop_lsuCoOp[3 : 0] <<< preShiftSize);
  assign stage1Out_payload_lsCtrlBundle_normalMemOp = ((stage1Out_payload_lsCtrlBundle_load || stage1Out_payload_lsCtrlBundle_store) && (! io_ctrl_stall));
  assign switch_LSU_l94 = io_input_payload_uop_lsuCoOp[3 : 0];
  always @(*) begin
    if((switch_LSU_l94 == LSUSizeOp_byte_1)) begin
        stage1Out_payload_lsCtrlBundle_size = 3'b000;
    end else if((switch_LSU_l94 == LSUSizeOp_halfword)) begin
        stage1Out_payload_lsCtrlBundle_size = {2'd0, _zz_stage1Out_payload_lsCtrlBundle_size};
    end else if((switch_LSU_l94 == LSUSizeOp_word)) begin
        stage1Out_payload_lsCtrlBundle_size = {1'd0, _zz_stage1Out_payload_lsCtrlBundle_size_1};
    end else begin
        stage1Out_payload_lsCtrlBundle_size = {1'd0, _zz_stage1Out_payload_lsCtrlBundle_size_2};
    end
  end

  assign stage1Out_payload_checkTLBException = (stage1Out_payload_lsCtrlBundle_normalMemOp || ((io_input_payload_uop_lsuOp == LSUOp_cacop) && (io_input_payload_uop_lsuCoOp == _zz_stage1Out_payload_checkTLBException)));
  assign stage1Out_payload_lsException = (! io_input_payload_exceptionInfo_exception);
  assign transferRAddr = {{transferRAddrHi,transferRAddrMid},transferRAddrLo};
  assign transferWAddr = {{transferWAddrHi,transferWAddrMid},transferWAddrLo};
  assign transferWriteBufferIdx = 3'b000;
  always @(*) begin
    mergedWrite[7 : 0] = ((transferLSMask[0] && missingEntry_store) ? transferWData[7 : 0] : io_axi_rdata[7 : 0]);
    mergedWrite[15 : 8] = ((transferLSMask[1] && missingEntry_store) ? transferWData[15 : 8] : io_axi_rdata[15 : 8]);
    mergedWrite[23 : 16] = ((transferLSMask[2] && missingEntry_store) ? transferWData[23 : 16] : io_axi_rdata[23 : 16]);
    mergedWrite[31 : 24] = ((transferLSMask[3] && missingEntry_store) ? transferWData[31 : 24] : io_axi_rdata[31 : 24]);
  end

  assign portAddr0 = (rollingBack ? latestWrite_index : _zz_portAddr0[10 : 2]);
  assign portWData0 = latestWrite_prevData;
  assign portWMask0 = 4'b1111;
  assign _zz_portRen0_0 = {stage1Out_ready,{stage1Out_ready,{stage1Out_ready,stage1Out_ready}}};
  assign portRen0_0 = (_zz_portRen0_0[0] || portWen0_0);
  assign portRen0_1 = (_zz_portRen0_0[1] || portWen0_1);
  assign portRen0_2 = (_zz_portRen0_0[2] || portWen0_2);
  assign portRen0_3 = (_zz_portRen0_0[3] || portWen0_3);
  assign _zz_portWen0_0 = {rollingBack,{rollingBack,{rollingBack,rollingBack}}};
  assign _zz_portWen0_0_1 = (! latestWrite_miss);
  assign _zz_portWen0_0_2 = {_zz_portWen0_0_1,{_zz_portWen0_0_1,{_zz_portWen0_0_1,_zz_portWen0_0_1}}};
  assign portWen0_0 = ((latestWrite_waySelect[0] && _zz_portWen0_0[0]) && _zz_portWen0_0_2[0]);
  assign portWen0_1 = ((latestWrite_waySelect[1] && _zz_portWen0_0[1]) && _zz_portWen0_0_2[1]);
  assign portWen0_2 = ((latestWrite_waySelect[2] && _zz_portWen0_0[2]) && _zz_portWen0_0_2[2]);
  assign portWen0_3 = ((latestWrite_waySelect[3] && _zz_portWen0_0[3]) && _zz_portWen0_0_2[3]);
  assign portAddr1 = (refilling ? ((io_axi_rready || io_axi_arvalid) ? _zz_portAddr1[10 : 2] : _zz_portAddr1_1[10 : 2]) : stage2In_payload_vaddr[10 : 2]);
  assign portWData1 = (refilling ? (writeBufferUpdate ? mergedWrite : io_axi_rdata) : stage2In_payload_storeData);
  assign portWMask1 = (refilling ? 4'b1111 : realLSMask);
  assign _zz_portRen1_0 = (io_axi_wready || io_axi_awvalid);
  assign _zz_portRen1_0_1 = {_zz_portRen1_0,{_zz_portRen1_0,{_zz_portRen1_0,_zz_portRen1_0}}};
  assign portRen1_0 = (_zz_portRen1_0_1[0] || portWen1_0);
  assign portRen1_1 = (_zz_portRen1_0_1[1] || portWen1_1);
  assign portRen1_2 = (_zz_portRen1_0_1[2] || portWen1_2);
  assign portRen1_3 = (_zz_portRen1_0_1[3] || portWen1_3);
  assign _zz_portWen1_1 = transferWaySelect[1];
  assign _zz_portWen1_2 = transferWaySelect[2];
  assign _zz_portWen1_3 = transferWaySelect[3];
  assign _zz_portWen1_0 = (io_axi_rvalid && io_axi_rready);
  assign _zz_portWen1_0_1 = {_zz_portWen1_0,{_zz_portWen1_0,{_zz_portWen1_0,_zz_portWen1_0}}};
  assign _zz_portWen1_1_1 = hit[1];
  assign _zz_portWen1_2_1 = hit[2];
  assign _zz_portWen1_3_1 = hit[3];
  assign _zz_portWen1_0_2 = (! miss);
  assign _zz_portWen1_0_3 = {_zz_portWen1_0_2,{_zz_portWen1_0_2,{_zz_portWen1_0_2,_zz_portWen1_0_2}}};
  assign _zz_portWen1_0_4 = {writeBufferAppend,{writeBufferAppend,{writeBufferAppend,writeBufferAppend}}};
  assign _zz_portWen1_0_5 = (! io_flush);
  assign _zz_portWen1_0_6 = {_zz_portWen1_0_5,{_zz_portWen1_0_5,{_zz_portWen1_0_5,_zz_portWen1_0_5}}};
  assign portWen1_0 = ((transferWaySelect[0] && _zz_portWen1_0_1[0]) || (((hit[0] && _zz_portWen1_0_3[0]) && _zz_portWen1_0_4[0]) && _zz_portWen1_0_6[0]));
  assign portWen1_1 = ((_zz_portWen1_1 && _zz_portWen1_0_1[1]) || (((_zz_portWen1_1_1 && _zz_portWen1_0_3[1]) && _zz_portWen1_0_4[1]) && _zz_portWen1_0_6[1]));
  assign portWen1_2 = ((_zz_portWen1_2 && _zz_portWen1_0_1[2]) || (((_zz_portWen1_2_1 && _zz_portWen1_0_3[2]) && _zz_portWen1_0_4[2]) && _zz_portWen1_0_6[2]));
  assign portWen1_3 = ((_zz_portWen1_3 && _zz_portWen1_0_1[3]) || (((_zz_portWen1_3_1 && _zz_portWen1_0_3[3]) && _zz_portWen1_0_4[3]) && _zz_portWen1_0_6[3]));
  always @(*) begin
    portRData0_0[7 : 0] = (portWMask1Bypass_0[0] ? portWData1Bypass_0[7 : 0] : portRData0Raw_0[7 : 0]);
    portRData0_0[15 : 8] = (portWMask1Bypass_0[1] ? portWData1Bypass_0[15 : 8] : portRData0Raw_0[15 : 8]);
    portRData0_0[23 : 16] = (portWMask1Bypass_0[2] ? portWData1Bypass_0[23 : 16] : portRData0Raw_0[23 : 16]);
    portRData0_0[31 : 24] = (portWMask1Bypass_0[3] ? portWData1Bypass_0[31 : 24] : portRData0Raw_0[31 : 24]);
  end

  assign when_LSU_l174 = (portWen1_0 && (portAddr0 == portAddr1));
  always @(*) begin
    portRData0_1[7 : 0] = (portWMask1Bypass_1[0] ? portWData1Bypass_1[7 : 0] : portRData0Raw_1[7 : 0]);
    portRData0_1[15 : 8] = (portWMask1Bypass_1[1] ? portWData1Bypass_1[15 : 8] : portRData0Raw_1[15 : 8]);
    portRData0_1[23 : 16] = (portWMask1Bypass_1[2] ? portWData1Bypass_1[23 : 16] : portRData0Raw_1[23 : 16]);
    portRData0_1[31 : 24] = (portWMask1Bypass_1[3] ? portWData1Bypass_1[31 : 24] : portRData0Raw_1[31 : 24]);
  end

  assign when_LSU_l174_1 = (portWen1_1 && (portAddr0 == portAddr1));
  always @(*) begin
    portRData0_2[7 : 0] = (portWMask1Bypass_2[0] ? portWData1Bypass_2[7 : 0] : portRData0Raw_2[7 : 0]);
    portRData0_2[15 : 8] = (portWMask1Bypass_2[1] ? portWData1Bypass_2[15 : 8] : portRData0Raw_2[15 : 8]);
    portRData0_2[23 : 16] = (portWMask1Bypass_2[2] ? portWData1Bypass_2[23 : 16] : portRData0Raw_2[23 : 16]);
    portRData0_2[31 : 24] = (portWMask1Bypass_2[3] ? portWData1Bypass_2[31 : 24] : portRData0Raw_2[31 : 24]);
  end

  assign when_LSU_l174_2 = (portWen1_2 && (portAddr0 == portAddr1));
  always @(*) begin
    portRData0_3[7 : 0] = (portWMask1Bypass_3[0] ? portWData1Bypass_3[7 : 0] : portRData0Raw_3[7 : 0]);
    portRData0_3[15 : 8] = (portWMask1Bypass_3[1] ? portWData1Bypass_3[15 : 8] : portRData0Raw_3[15 : 8]);
    portRData0_3[23 : 16] = (portWMask1Bypass_3[2] ? portWData1Bypass_3[23 : 16] : portRData0Raw_3[23 : 16]);
    portRData0_3[31 : 24] = (portWMask1Bypass_3[3] ? portWData1Bypass_3[31 : 24] : portRData0Raw_3[31 : 24]);
  end

  assign when_LSU_l174_3 = (portWen1_3 && (portAddr0 == portAddr1));
  always @(*) begin
    stage1Out_payload_wayValid[0] = _zz_stage1Out_payload_wayValid;
    stage1Out_payload_wayValid[1] = _zz_stage1Out_payload_wayValid_3;
    stage1Out_payload_wayValid[2] = _zz_stage1Out_payload_wayValid_6;
    stage1Out_payload_wayValid[3] = _zz_stage1Out_payload_wayValid_9;
  end

  always @(*) begin
    stage1Out_payload_wayDirty[0] = _zz_stage1Out_payload_wayDirty;
    stage1Out_payload_wayDirty[1] = _zz_stage1Out_payload_wayDirty_3;
    stage1Out_payload_wayDirty[2] = _zz_stage1Out_payload_wayDirty_6;
    stage1Out_payload_wayDirty[3] = _zz_stage1Out_payload_wayDirty_9;
  end

  assign dataRead_0 = portRData0_0;
  assign portRData0Raw_0 = data_0_portA_rdData;
  assign portRData1_0 = data_0_portB_rdData;
  assign stage1Out_fire = (stage1Out_valid && stage1Out_ready);
  assign tagRead_0 = tag_0_rd_data;
  always @(*) begin
    hit[0] = ((stage2In_payload_wayValid[0] && (tagRead_0 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_vaddr[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit));
    hit[1] = ((stage2In_payload_wayValid[1] && (tagRead_1 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_vaddr[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit_2));
    hit[2] = ((stage2In_payload_wayValid[2] && (tagRead_2 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_vaddr[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit_4));
    hit[3] = ((stage2In_payload_wayValid[3] && (tagRead_3 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_vaddr[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit_6));
  end

  assign dataRead_1 = portRData0_1;
  assign portRData0Raw_1 = data_1_portA_rdData;
  assign portRData1_1 = data_1_portB_rdData;
  assign tagRead_1 = tag_1_rd_data;
  assign dataRead_2 = portRData0_2;
  assign portRData0Raw_2 = data_2_portA_rdData;
  assign portRData1_2 = data_2_portB_rdData;
  assign tagRead_2 = tag_2_rd_data;
  assign dataRead_3 = portRData0_3;
  assign portRData0Raw_3 = data_3_portA_rdData;
  assign portRData1_3 = data_3_portB_rdData;
  assign tagRead_3 = tag_3_rd_data;
  assign miss = ((stage2In_valid && stage2In_payload_lsCtrlBundle_normalMemOp) && (! ((|hit) || exceptionInfo_exception)));
  assign _zz_exceptionInfo_exception = (stage2In_payload_exceptionInfo_exception || (! stage2In_payload_checkTLBException));
  assign exceptionInfo_exception = (_zz_exceptionInfo_exception ? stage1Out_payload_exceptionInfo_exception : exceptionInfo2_exception);
  assign exceptionInfo_eCode = (_zz_exceptionInfo_exception ? stage1Out_payload_exceptionInfo_eCode : exceptionInfo2_eCode);
  assign exceptionInfo_eSubCode = (_zz_exceptionInfo_exception ? stage1Out_payload_exceptionInfo_eSubCode : exceptionInfo2_eSubCode);
  assign noStructuralHazard = (((! axiLoad) && ((! miss) || missBufferAvail)) && ((! stage2In_payload_lsCtrlBundle_store) || writeBufferAvail));
  always @(*) begin
    axiFinish = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
      end
      axiCtrl_enumDef_readReq : begin
      end
      axiCtrl_enumDef_readFirst : begin
      end
      axiCtrl_enumDef_read : begin
        if(when_LSU_l510) begin
          if(io_axi_rlast) begin
            axiFinish = 1'b1;
          end
        end
      end
      axiCtrl_enumDef_writeReq : begin
      end
      axiCtrl_enumDef_write : begin
        if(when_LSU_l539) begin
          if(io_axi_wlast) begin
            if(transferUncached) begin
              axiFinish = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign stage2In_ready = (noStructuralHazard || io_flush);
  assign when_LSU_l203 = (((stage1Out_payload_lsCtrlBundle_load || stage1Out_payload_lsCtrlBundle_store) && ((io_input_payload_uop_lsuCoOp[3 : 0] == LSUSizeOp_word) && (|address[1 : 0]))) || ((io_input_payload_uop_lsuCoOp[3 : 0] == LSUSizeOp_halfword) && address[0]));
  always @(*) begin
    if(when_LSU_l203) begin
      exceptionInfo1_exception = 1'b1;
    end else begin
      exceptionInfo1_exception = 1'b0;
    end
  end

  always @(*) begin
    if(when_LSU_l203) begin
      exceptionInfo1_eCode = {2'd0, _zz_exceptionInfo1_eCode};
    end else begin
      exceptionInfo1_eCode = {2'd0, _zz_exceptionInfo1_eCode_1};
    end
  end

  always @(*) begin
    if(when_LSU_l203) begin
      exceptionInfo1_eSubCode = 1'b0;
    end else begin
      exceptionInfo1_eSubCode = 1'b0;
    end
  end

  assign when_LSU_l213 = (! stage2In_payload_tlb_pageInfo_v);
  always @(*) begin
    if(stage2In_payload_tlb_hit) begin
      if(when_LSU_l213) begin
        exceptionInfo2_exception = 1'b1;
      end else begin
        if(when_LSU_l217) begin
          exceptionInfo2_exception = 1'b1;
        end else begin
          if(when_LSU_l221) begin
            exceptionInfo2_exception = 1'b1;
          end else begin
            exceptionInfo2_exception = 1'b0;
          end
        end
      end
    end else begin
      exceptionInfo2_exception = 1'b1;
    end
  end

  always @(*) begin
    if(stage2In_payload_tlb_hit) begin
      if(when_LSU_l213) begin
        exceptionInfo2_eCode = (stage2In_payload_lsCtrlBundle_load ? _zz_exceptionInfo2_eCode : _zz_exceptionInfo2_eCode_2);
      end else begin
        if(when_LSU_l217) begin
          exceptionInfo2_eCode = {3'd0, _zz_exceptionInfo2_eCode_4};
        end else begin
          if(when_LSU_l221) begin
            exceptionInfo2_eCode = {3'd0, _zz_exceptionInfo2_eCode_5};
          end else begin
            exceptionInfo2_eCode = {3'd0, _zz_exceptionInfo2_eCode_6};
          end
        end
      end
    end else begin
      exceptionInfo2_eCode = 6'h3f;
    end
  end

  always @(*) begin
    if(stage2In_payload_tlb_hit) begin
      if(when_LSU_l213) begin
        exceptionInfo2_eSubCode = (stage2In_payload_lsCtrlBundle_load ? 1'b0 : 1'b0);
      end else begin
        if(when_LSU_l217) begin
          exceptionInfo2_eSubCode = 1'b0;
        end else begin
          if(when_LSU_l221) begin
            exceptionInfo2_eSubCode = 1'b0;
          end else begin
            exceptionInfo2_eSubCode = 1'b0;
          end
        end
      end
    end else begin
      exceptionInfo2_eSubCode = 1'b0;
    end
  end

  assign when_LSU_l217 = (stage2In_payload_tlb_pageInfo_plv < _zz_when_LSU_l217);
  assign when_LSU_l221 = (stage2In_payload_lsCtrlBundle_store && (! stage2In_payload_tlb_pageInfo_d));
  assign scMatchHit = ((stage2In_payload_lsCtrlBundle_sc && ({stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_vaddr[11 : 0]} == io_llBitComm_actualAddr)) && _zz_scMatchHit);
  assign scMatchAXI = ((missingEntry_sc && (transferRAddr == io_llBitComm_actualAddr)) && _zz_scMatchHit);
  assign scResHit = {31'h00000000,scMatchHit};
  assign scResAXI = {31'h00000000,scMatchAXI};
  assign realLSMask = ((stage2In_payload_lsCtrlBundle_sc && (! scMatchHit)) ? 4'b0000 : stage2In_payload_lsCtrlBundle_lsMask);
  assign io_llBitComm_toUpdateAddr = {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_vaddr[11 : 0]};
  assign io_llBitComm_wen = (stage2In_payload_lsCtrlBundle_ll && stage2In_valid);
  assign _zz_writeBufferHeadNext = 4'b0000;
  assign _zz_writeBufferHeadNext_1 = 4'b0001;
  assign _zz_writeBufferHeadNext_2 = 4'b0001;
  assign _zz_writeBufferHeadNext_3 = 4'b0010;
  assign _zz_writeBufferHeadNext_4 = 4'b0001;
  assign _zz_writeBufferHeadNext_5 = 4'b0010;
  assign _zz_writeBufferHeadNext_6 = 4'b0010;
  assign _zz_writeBufferHeadNext_7 = 4'b0011;
  assign writeBufferHeadNext = (writeBufferHead + _zz_writeBufferHeadNext_8);
  assign _zz_writeBufferAvail = _zz__zz_writeBufferAvail;
  assign _zz_1 = ({7'd0,1'b1} <<< writeBufferTail);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = _zz_1[4];
  assign _zz_7 = _zz_1[5];
  assign _zz_8 = _zz_1[6];
  assign _zz_9 = _zz_1[7];
  assign latestWrite_robIdx = _zz_latestWrite_robIdx;
  assign latestWrite_waySelect = _zz_latestWrite_waySelect;
  assign latestWrite_prevData = _zz_latestWrite_prevData;
  assign latestWrite_prevDirty = _zz_latestWrite_prevDirty;
  assign latestWrite_index = _zz_latestWrite_index;
  assign latestWrite_miss = _zz_latestWrite_miss;
  assign latestWrite_valid = _zz_writeBufferAvail;
  assign writeBufferAvail = (! _zz_writeBufferAvail);
  always @(*) begin
    _zz_writeBufferRetireMask[0] = ((writeBuffer_0_robIdx == io_retireComm_robIdx_0) && io_retireComm_allowRetire_0);
    _zz_writeBufferRetireMask[1] = ((writeBuffer_0_robIdx == io_retireComm_robIdx_1) && io_retireComm_allowRetire_1);
  end

  always @(*) begin
    writeBufferRetireMask[0] = ((|_zz_writeBufferRetireMask) && writeBuffer_0_valid);
    writeBufferRetireMask[1] = ((|_zz_writeBufferRetireMask_1) && writeBuffer_1_valid);
    writeBufferRetireMask[2] = ((|_zz_writeBufferRetireMask_2) && writeBuffer_2_valid);
    writeBufferRetireMask[3] = ((|_zz_writeBufferRetireMask_3) && writeBuffer_3_valid);
    writeBufferRetireMask[4] = ((|_zz_writeBufferRetireMask_4) && writeBuffer_4_valid);
    writeBufferRetireMask[5] = ((|_zz_writeBufferRetireMask_5) && writeBuffer_5_valid);
    writeBufferRetireMask[6] = ((|_zz_writeBufferRetireMask_6) && writeBuffer_6_valid);
    writeBufferRetireMask[7] = ((|_zz_writeBufferRetireMask_7) && writeBuffer_7_valid);
  end

  always @(*) begin
    _zz_writeBufferRetireMask_1[0] = ((writeBuffer_1_robIdx == io_retireComm_robIdx_0) && io_retireComm_allowRetire_0);
    _zz_writeBufferRetireMask_1[1] = ((writeBuffer_1_robIdx == io_retireComm_robIdx_1) && io_retireComm_allowRetire_1);
  end

  always @(*) begin
    _zz_writeBufferRetireMask_2[0] = ((writeBuffer_2_robIdx == io_retireComm_robIdx_0) && io_retireComm_allowRetire_0);
    _zz_writeBufferRetireMask_2[1] = ((writeBuffer_2_robIdx == io_retireComm_robIdx_1) && io_retireComm_allowRetire_1);
  end

  always @(*) begin
    _zz_writeBufferRetireMask_3[0] = ((writeBuffer_3_robIdx == io_retireComm_robIdx_0) && io_retireComm_allowRetire_0);
    _zz_writeBufferRetireMask_3[1] = ((writeBuffer_3_robIdx == io_retireComm_robIdx_1) && io_retireComm_allowRetire_1);
  end

  always @(*) begin
    _zz_writeBufferRetireMask_4[0] = ((writeBuffer_4_robIdx == io_retireComm_robIdx_0) && io_retireComm_allowRetire_0);
    _zz_writeBufferRetireMask_4[1] = ((writeBuffer_4_robIdx == io_retireComm_robIdx_1) && io_retireComm_allowRetire_1);
  end

  always @(*) begin
    _zz_writeBufferRetireMask_5[0] = ((writeBuffer_5_robIdx == io_retireComm_robIdx_0) && io_retireComm_allowRetire_0);
    _zz_writeBufferRetireMask_5[1] = ((writeBuffer_5_robIdx == io_retireComm_robIdx_1) && io_retireComm_allowRetire_1);
  end

  always @(*) begin
    _zz_writeBufferRetireMask_6[0] = ((writeBuffer_6_robIdx == io_retireComm_robIdx_0) && io_retireComm_allowRetire_0);
    _zz_writeBufferRetireMask_6[1] = ((writeBuffer_6_robIdx == io_retireComm_robIdx_1) && io_retireComm_allowRetire_1);
  end

  always @(*) begin
    _zz_writeBufferRetireMask_7[0] = ((writeBuffer_7_robIdx == io_retireComm_robIdx_0) && io_retireComm_allowRetire_0);
    _zz_writeBufferRetireMask_7[1] = ((writeBuffer_7_robIdx == io_retireComm_robIdx_1) && io_retireComm_allowRetire_1);
  end

  assign writeBufferAppend = (((((stage2In_payload_lsCtrlBundle_store && (stage2In_payload_tlb_pageInfo_mat == _zz_writeBufferAppend)) && stage2In_valid) && (! exceptionInfo_exception)) && noStructuralHazard) && (! cacopActive));
  assign when_LSU_l267 = (writeBufferAppend && (! io_flush));
  assign _zz_writeBuffer_0_waySelect = (miss ? wayToReplace : hit);
  assign _zz_io_output_payload_data = (_zz_portWen1_1_1 || _zz_portWen1_3_1);
  assign _zz_io_output_payload_data_1 = (_zz_portWen1_2_1 || _zz_portWen1_3_1);
  assign _zz_io_output_payload_data_2 = {_zz_io_output_payload_data_1,_zz_io_output_payload_data};
  assign _zz_writeBuffer_0_prevData = _zz__zz_writeBuffer_0_prevData;
  assign _zz_missBuffer_0_writeBack = wayDirty[0];
  assign _zz_missBuffer_0_writeBack_1 = wayDirty[1];
  assign _zz_missBuffer_0_writeBack_2 = wayDirty[2];
  assign _zz_missBuffer_0_writeBack_3 = wayDirty[3];
  assign _zz_writeBuffer_0_prevDirty = (miss ? 1'b0 : _zz__zz_writeBuffer_0_prevDirty);
  assign _zz_writeBuffer_0_index = stage2In_payload_vaddr[10 : 2];
  assign _zz_10 = ({7'd0,1'b1} <<< missingEntry_writeBufferIdx);
  assign _zz_11 = _zz_10[0];
  assign _zz_12 = _zz_10[1];
  assign _zz_13 = _zz_10[2];
  assign _zz_14 = _zz_10[3];
  assign _zz_15 = _zz_10[4];
  assign _zz_16 = _zz_10[5];
  assign _zz_17 = _zz_10[6];
  assign _zz_18 = _zz_10[7];
  assign missingEntry_robIdx = missBuffer_0_robIdx;
  assign missingEntry_prd = missBuffer_0_prd;
  assign missingEntry_branchResult_targetPC = missBuffer_0_branchResult_targetPC;
  assign missingEntry_branchResult_branchResult = missBuffer_0_branchResult_branchResult;
  assign missingEntry_branchResult_predictFail = missBuffer_0_branchResult_predictFail;
  assign missingEntry_exceptionInfo_exception = missBuffer_0_exceptionInfo_exception;
  assign missingEntry_exceptionInfo_eCode = missBuffer_0_exceptionInfo_eCode;
  assign missingEntry_exceptionInfo_eSubCode = missBuffer_0_exceptionInfo_eSubCode;
  assign missingEntry_uncached = missBuffer_0_uncached;
  assign missingEntry_load = missBuffer_0_load;
  assign missingEntry_store = missBuffer_0_store;
  assign missingEntry_signed = missBuffer_0_signed;
  assign missingEntry_ll = missBuffer_0_ll;
  assign missingEntry_sc = missBuffer_0_sc;
  assign missingEntry_writeBufferIdx = missBuffer_0_writeBufferIdx;
  assign missingEntry_waySelect = missBuffer_0_waySelect;
  assign missingEntry_writeBack = missBuffer_0_writeBack;
  assign missingEntry_storeData = missBuffer_0_storeData;
  assign missingEntry_lsMask = missBuffer_0_lsMask;
  assign missingEntry_size = missBuffer_0_size;
  assign missingEntry_vaddr = missBuffer_0_vaddr;
  assign missingEntry_paddr = missBuffer_0_paddr;
  assign missingEntry_prevPaddr = missBuffer_0_prevPaddr;
  assign missingEntry_valid = missBuffer_0_valid;
  assign _zz_19 = _zz__zz_19[0];
  assign missBufferAvail = (! missBuffer_0_valid);
  assign when_LSU_l292 = ((miss && stage2In_ready) && (! io_flush));
  assign _zz_missBuffer_0_writeBack_4 = wayToReplace[3];
  assign _zz_missBuffer_0_writeBack_5 = (wayToReplace[1] || _zz_missBuffer_0_writeBack_4);
  assign _zz_missBuffer_0_writeBack_6 = (wayToReplace[2] || _zz_missBuffer_0_writeBack_4);
  assign _zz_missBuffer_0_writeBack_7 = {_zz_missBuffer_0_writeBack_6,_zz_missBuffer_0_writeBack_5};
  always @(*) begin
    sameBlockMask[0] = ((missBuffer_0_valid && (! missBuffer_0_uncached)) && (missBuffer_0_vaddr[10 : 6] == address[10 : 6]));
    sameBlockMask[1] = ((miss && (! (stage2In_payload_tlb_pageInfo_mat == 2'b00))) && (stage2In_payload_vaddr[10 : 6] == address[10 : 6]));
  end

  assign sameBlock = ((|sameBlockMask) && io_input_valid);
  assign stall = ((io_ctrl_stall || sameBlock) || rollingBack);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_LSU_l335 = ((io_output_fire && (axiLoad ? (! transferUncached) : (stage2In_payload_lsCtrlBundle_normalMemOp && (stage2In_payload_tlb_pageInfo_mat == _zz_when_LSU_l335)))) && (! exceptionInfo_exception));
  assign _zz_20 = ({31'd0,1'b1} <<< (axiLoad ? missingEntry_vaddr[10 : 6] : stage2In_payload_vaddr[10 : 6]));
  assign _zz_21 = _zz_20[0];
  assign _zz_22 = _zz_20[1];
  assign _zz_23 = _zz_20[2];
  assign _zz_24 = _zz_20[3];
  assign _zz_25 = _zz_20[4];
  assign _zz_26 = _zz_20[5];
  assign _zz_27 = _zz_20[6];
  assign _zz_28 = _zz_20[7];
  assign _zz_29 = _zz_20[8];
  assign _zz_30 = _zz_20[9];
  assign _zz_31 = _zz_20[10];
  assign _zz_32 = _zz_20[11];
  assign _zz_33 = _zz_20[12];
  assign _zz_34 = _zz_20[13];
  assign _zz_35 = _zz_20[14];
  assign _zz_36 = _zz_20[15];
  assign _zz_37 = _zz_20[16];
  assign _zz_38 = _zz_20[17];
  assign _zz_39 = _zz_20[18];
  assign _zz_40 = _zz_20[19];
  assign _zz_41 = _zz_20[20];
  assign _zz_42 = _zz_20[21];
  assign _zz_43 = _zz_20[22];
  assign _zz_44 = _zz_20[23];
  assign _zz_45 = _zz_20[24];
  assign _zz_46 = _zz_20[25];
  assign _zz_47 = _zz_20[26];
  assign _zz_48 = _zz_20[27];
  assign _zz_49 = _zz_20[28];
  assign _zz_50 = _zz_20[29];
  assign _zz_51 = _zz_20[30];
  assign _zz_52 = _zz_20[31];
  assign _zz_lruBit_0_0 = (axiLoad ? (|transferWaySelect[3 : 2]) : (|hit[3 : 2]));
  assign _zz_lruBit_0_1 = (axiLoad ? (|transferWaySelect[1 : 1]) : (|hit[1 : 1]));
  assign _zz_lruBit_0_2 = (axiLoad ? (|transferWaySelect[3 : 3]) : (|hit[3 : 3]));
  assign dirtyUpdate = ((io_output_fire && (axiLoad ? ((! transferUncached) && missingEntry_store) : (stage2In_payload_lsCtrlBundle_store && (stage2In_payload_tlb_pageInfo_mat == _zz_dirtyUpdate)))) && (! exceptionInfo_exception));
  assign when_LSU_l341 = (axiLoad ? transferWaySelect[0] : hit[0]);
  assign _zz_53 = ({31'd0,1'b1} <<< (axiLoad ? _zz__zz_53[10 : 6] : stage2In_payload_vaddr[10 : 6]));
  assign when_LSU_l341_1 = (axiLoad ? transferWaySelect[1] : hit[1]);
  assign _zz_54 = ({31'd0,1'b1} <<< (axiLoad ? _zz__zz_54[10 : 6] : stage2In_payload_vaddr[10 : 6]));
  assign when_LSU_l341_2 = (axiLoad ? transferWaySelect[2] : hit[2]);
  assign _zz_55 = ({31'd0,1'b1} <<< (axiLoad ? _zz__zz_55[10 : 6] : stage2In_payload_vaddr[10 : 6]));
  assign when_LSU_l341_3 = (axiLoad ? transferWaySelect[3] : hit[3]);
  assign _zz_56 = ({31'd0,1'b1} <<< (axiLoad ? _zz__zz_56[10 : 6] : stage2In_payload_vaddr[10 : 6]));
  assign when_LSU_l348 = latestWrite_waySelect[0];
  assign _zz_57 = ({31'd0,1'b1} <<< latestWrite_index[8 : 4]);
  assign when_LSU_l348_1 = latestWrite_waySelect[1];
  assign _zz_58 = ({31'd0,1'b1} <<< latestWrite_index[8 : 4]);
  assign when_LSU_l348_2 = latestWrite_waySelect[2];
  assign _zz_59 = ({31'd0,1'b1} <<< latestWrite_index[8 : 4]);
  assign when_LSU_l348_3 = latestWrite_waySelect[3];
  assign _zz_60 = ({31'd0,1'b1} <<< latestWrite_index[8 : 4]);
  assign wayDirty = (stage2In_payload_wayDirty | wayDirtyBypass);
  assign when_LSU_l357 = (dirtyUpdate && ((axiLoad ? _zz_when_LSU_l357[10 : 6] : stage2In_payload_vaddr[10 : 6]) == _zz_when_LSU_l357_1[10 : 6]));
  assign io_axi_arid = {3'd0, _zz_io_axi_arid};
  assign io_axi_araddr = (transferUncached ? transferRAddr : {transferRAddr[31 : 2],2'b00});
  assign io_axi_arlen = (transferUncached ? 8'h00 : _zz_io_axi_arlen);
  assign io_axi_arsize = (transferUncached ? missingEntry_size : _zz_io_axi_arsize);
  assign io_axi_arburst = (transferUncached ? 2'b01 : 2'b10);
  assign io_axi_arlock = 2'b00;
  assign io_axi_arcache = 4'b0000;
  assign io_axi_arprot = 3'b000;
  always @(*) begin
    io_axi_arvalid = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
        io_axi_arvalid = 1'b0;
      end
      axiCtrl_enumDef_readReq : begin
        io_axi_arvalid = 1'b1;
      end
      axiCtrl_enumDef_readFirst : begin
        io_axi_arvalid = 1'b0;
      end
      axiCtrl_enumDef_read : begin
        io_axi_arvalid = 1'b0;
      end
      axiCtrl_enumDef_writeReq : begin
        io_axi_arvalid = 1'b0;
      end
      axiCtrl_enumDef_write : begin
        io_axi_arvalid = 1'b0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_rready = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
        io_axi_rready = 1'b0;
      end
      axiCtrl_enumDef_readReq : begin
        io_axi_rready = 1'b0;
      end
      axiCtrl_enumDef_readFirst : begin
        io_axi_rready = 1'b1;
      end
      axiCtrl_enumDef_read : begin
        io_axi_rready = 1'b1;
      end
      axiCtrl_enumDef_writeReq : begin
        io_axi_rready = 1'b0;
      end
      axiCtrl_enumDef_write : begin
        io_axi_rready = 1'b0;
      end
      default : begin
      end
    endcase
  end

  assign io_axi_awid = {3'd0, _zz_io_axi_awid};
  assign io_axi_awaddr = transferWAddr;
  assign io_axi_awlen = {4'd0, _zz_io_axi_awlen};
  assign io_axi_awsize = (transferUncached ? missingEntry_size : _zz_io_axi_awsize);
  assign io_axi_awburst = {1'd0, _zz_io_axi_awburst};
  assign io_axi_awlock = 2'b00;
  assign io_axi_awcache = 4'b0000;
  assign io_axi_awprot = 3'b000;
  always @(*) begin
    io_axi_awvalid = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
        io_axi_awvalid = 1'b0;
      end
      axiCtrl_enumDef_readReq : begin
        io_axi_awvalid = 1'b0;
      end
      axiCtrl_enumDef_readFirst : begin
        io_axi_awvalid = 1'b0;
      end
      axiCtrl_enumDef_read : begin
        io_axi_awvalid = 1'b0;
      end
      axiCtrl_enumDef_writeReq : begin
        io_axi_awvalid = 1'b1;
      end
      axiCtrl_enumDef_write : begin
        io_axi_awvalid = 1'b0;
      end
      default : begin
      end
    endcase
  end

  assign io_axi_wid = {3'd0, _zz_io_axi_wid};
  assign _zz_io_axi_wdata = (_zz_portWen1_1 || _zz_portWen1_3);
  assign _zz_io_axi_wdata_1 = (_zz_portWen1_2 || _zz_portWen1_3);
  assign io_axi_wdata = (transferUncached ? transferWData : _zz_io_axi_wdata_2);
  assign io_axi_wstrb = (transferUncached ? transferLSMask : 4'b1111);
  assign io_axi_wlast = ((&transferWAddrMid) || transferUncached);
  always @(*) begin
    io_axi_wvalid = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
        io_axi_wvalid = 1'b0;
      end
      axiCtrl_enumDef_readReq : begin
        io_axi_wvalid = 1'b0;
      end
      axiCtrl_enumDef_readFirst : begin
        io_axi_wvalid = 1'b0;
      end
      axiCtrl_enumDef_read : begin
        io_axi_wvalid = 1'b0;
      end
      axiCtrl_enumDef_writeReq : begin
        io_axi_wvalid = 1'b0;
      end
      axiCtrl_enumDef_write : begin
        io_axi_wvalid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign io_axi_bready = 1'b1;
  always @(*) begin
    axiLoad = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
      end
      axiCtrl_enumDef_readReq : begin
      end
      axiCtrl_enumDef_readFirst : begin
        if(when_LSU_l496) begin
          axiLoad = 1'b1;
        end
      end
      axiCtrl_enumDef_read : begin
      end
      axiCtrl_enumDef_writeReq : begin
      end
      axiCtrl_enumDef_write : begin
        if(when_LSU_l539) begin
          if(io_axi_wlast) begin
            if(transferUncached) begin
              axiLoad = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    refilling = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
        refilling = 1'b0;
      end
      axiCtrl_enumDef_readReq : begin
        refilling = 1'b1;
      end
      axiCtrl_enumDef_readFirst : begin
        refilling = 1'b1;
      end
      axiCtrl_enumDef_read : begin
        refilling = 1'b1;
      end
      axiCtrl_enumDef_writeReq : begin
        refilling = 1'b1;
      end
      axiCtrl_enumDef_write : begin
        refilling = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    rollingBack = 1'b0;
    case(rollbackCtrl_stateReg)
      rollbackCtrl_enumDef_idle : begin
        rollingBack = 1'b0;
      end
      rollbackCtrl_enumDef_rollback : begin
        rollingBack = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    writeBufferUpdate = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
        writeBufferUpdate = 1'b0;
      end
      axiCtrl_enumDef_readReq : begin
        writeBufferUpdate = 1'b0;
      end
      axiCtrl_enumDef_readFirst : begin
        writeBufferUpdate = (missingEntry_store && (io_axi_rvalid && io_axi_rready));
      end
      axiCtrl_enumDef_read : begin
        writeBufferUpdate = 1'b0;
      end
      axiCtrl_enumDef_writeReq : begin
        writeBufferUpdate = 1'b0;
      end
      axiCtrl_enumDef_write : begin
        writeBufferUpdate = 1'b0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_missBufferAllowMask[0] = (missBuffer_0_robIdx == io_retireComm_robIdx_0);
    _zz_missBufferAllowMask[1] = ((missBuffer_0_robIdx == io_retireComm_robIdx_1) && (&_zz__zz_missBufferAllowMask[0 : 0]));
  end

  assign missBufferAllowMask[0] = (((|_zz_missBufferAllowMask) && missBuffer_0_valid) && (! io_flush));
  always @(*) begin
    _zz_missBufferPreAllowMask[0] = ((_zz__zz_missBufferPreAllowMask == writeBuffer_0_index) && writeBuffer_0_valid);
    _zz_missBufferPreAllowMask[1] = ((_zz__zz_missBufferPreAllowMask_2 == writeBuffer_1_index) && writeBuffer_1_valid);
    _zz_missBufferPreAllowMask[2] = ((_zz__zz_missBufferPreAllowMask_4 == writeBuffer_2_index) && writeBuffer_2_valid);
    _zz_missBufferPreAllowMask[3] = ((_zz__zz_missBufferPreAllowMask_6 == writeBuffer_3_index) && writeBuffer_3_valid);
    _zz_missBufferPreAllowMask[4] = ((_zz__zz_missBufferPreAllowMask_8 == writeBuffer_4_index) && writeBuffer_4_valid);
    _zz_missBufferPreAllowMask[5] = ((_zz__zz_missBufferPreAllowMask_10 == writeBuffer_5_index) && writeBuffer_5_valid);
    _zz_missBufferPreAllowMask[6] = ((_zz__zz_missBufferPreAllowMask_12 == writeBuffer_6_index) && writeBuffer_6_valid);
    _zz_missBufferPreAllowMask[7] = ((_zz__zz_missBufferPreAllowMask_14 == writeBuffer_7_index) && writeBuffer_7_valid);
  end

  assign missBufferPreAllowMask[0] = (((|_zz_missBufferPreAllowMask) && missBuffer_0_valid) && (! io_flush));
  assign cacopPAddr = (stage2In_payload_isHitInvalidate ? {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_vaddr[11 : 0]} : {{_zz_cacopPAddr,stage2In_payload_vaddr[10 : 6]},6'h00});
  assign axiCtrl_wantExit = 1'b0;
  always @(*) begin
    axiCtrl_wantStart = 1'b0;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
      end
      axiCtrl_enumDef_readReq : begin
      end
      axiCtrl_enumDef_readFirst : begin
      end
      axiCtrl_enumDef_read : begin
      end
      axiCtrl_enumDef_writeReq : begin
      end
      axiCtrl_enumDef_write : begin
      end
      default : begin
        axiCtrl_wantStart = 1'b1;
      end
    endcase
  end

  assign axiCtrl_wantKill = 1'b0;
  assign rollbackCtrl_wantExit = 1'b0;
  always @(*) begin
    rollbackCtrl_wantStart = 1'b0;
    case(rollbackCtrl_stateReg)
      rollbackCtrl_enumDef_idle : begin
      end
      rollbackCtrl_enumDef_rollback : begin
      end
      default : begin
        rollbackCtrl_wantStart = 1'b1;
      end
    endcase
  end

  assign rollbackCtrl_wantKill = 1'b0;
  always @(*) begin
    _zz_wayToReplace[0] = (! _zz__zz_wayToReplace);
    _zz_wayToReplace[1] = (! _zz__zz_wayToReplace_2);
  end

  always @(*) begin
    wayToReplace[0] = (&_zz_wayToReplace);
    wayToReplace[1] = (&_zz_wayToReplace_1);
    wayToReplace[2] = (&_zz_wayToReplace_2);
    wayToReplace[3] = (&_zz_wayToReplace_3);
  end

  always @(*) begin
    _zz_wayToReplace_1[0] = (! _zz__zz_wayToReplace_1_1);
    _zz_wayToReplace_1[1] = _zz__zz_wayToReplace_1_3;
  end

  always @(*) begin
    _zz_wayToReplace_2[0] = _zz__zz_wayToReplace_2_1;
    _zz_wayToReplace_2[1] = (! _zz__zz_wayToReplace_2_3);
  end

  always @(*) begin
    _zz_wayToReplace_3[0] = _zz__zz_wayToReplace_3_1;
    _zz_wayToReplace_3[1] = _zz__zz_wayToReplace_3_3;
  end

  assign _zz_dataShuffle_0 = (dataRead_0 >>> stage2In_payload_vaddr[5 : 0]);
  assign _zz_dataShuffle_0_1 = (_zz_dataShuffle_0[7] && stage2In_payload_lsCtrlBundle_signed);
  always @(*) begin
    case(stage2In_payload_lsCtrlBundle_size)
      3'b000 : begin
        dataShuffle_0 = {{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_1,{_zz_dataShuffle_0_3,_zz_dataShuffle_0_4}}}}}}}}}},_zz_dataShuffle_0[7 : 0]};
      end
      3'b001 : begin
        dataShuffle_0 = {{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_2,{_zz_dataShuffle_0_5,_zz_dataShuffle_0_6}}}}}}}}}},_zz_dataShuffle_0[15 : 0]};
      end
      3'b010 : begin
        dataShuffle_0 = _zz_dataShuffle_0;
      end
      default : begin
        dataShuffle_0 = _zz_dataShuffle_0;
      end
    endcase
  end

  assign _zz_dataShuffle_0_2 = (_zz_dataShuffle_0[15] && stage2In_payload_lsCtrlBundle_signed);
  assign _zz_dataShuffle_1 = (dataRead_1 >>> stage2In_payload_vaddr[5 : 0]);
  assign _zz_dataShuffle_1_1 = (_zz_dataShuffle_1[7] && stage2In_payload_lsCtrlBundle_signed);
  always @(*) begin
    case(stage2In_payload_lsCtrlBundle_size)
      3'b000 : begin
        dataShuffle_1 = {{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_1,{_zz_dataShuffle_1_3,_zz_dataShuffle_1_4}}}}}}}}}},_zz_dataShuffle_1[7 : 0]};
      end
      3'b001 : begin
        dataShuffle_1 = {{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_2,{_zz_dataShuffle_1_5,_zz_dataShuffle_1_6}}}}}}}}}},_zz_dataShuffle_1[15 : 0]};
      end
      3'b010 : begin
        dataShuffle_1 = _zz_dataShuffle_1;
      end
      default : begin
        dataShuffle_1 = _zz_dataShuffle_1;
      end
    endcase
  end

  assign _zz_dataShuffle_1_2 = (_zz_dataShuffle_1[15] && stage2In_payload_lsCtrlBundle_signed);
  assign _zz_dataShuffle_2 = (dataRead_2 >>> stage2In_payload_vaddr[5 : 0]);
  assign _zz_dataShuffle_2_1 = (_zz_dataShuffle_2[7] && stage2In_payload_lsCtrlBundle_signed);
  always @(*) begin
    case(stage2In_payload_lsCtrlBundle_size)
      3'b000 : begin
        dataShuffle_2 = {{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_1,{_zz_dataShuffle_2_3,_zz_dataShuffle_2_4}}}}}}}}}},_zz_dataShuffle_2[7 : 0]};
      end
      3'b001 : begin
        dataShuffle_2 = {{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_2,{_zz_dataShuffle_2_5,_zz_dataShuffle_2_6}}}}}}}}}},_zz_dataShuffle_2[15 : 0]};
      end
      3'b010 : begin
        dataShuffle_2 = _zz_dataShuffle_2;
      end
      default : begin
        dataShuffle_2 = _zz_dataShuffle_2;
      end
    endcase
  end

  assign _zz_dataShuffle_2_2 = (_zz_dataShuffle_2[15] && stage2In_payload_lsCtrlBundle_signed);
  assign _zz_dataShuffle_3 = (dataRead_3 >>> stage2In_payload_vaddr[5 : 0]);
  assign _zz_dataShuffle_3_1 = (_zz_dataShuffle_3[7] && stage2In_payload_lsCtrlBundle_signed);
  always @(*) begin
    case(stage2In_payload_lsCtrlBundle_size)
      3'b000 : begin
        dataShuffle_3 = {{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_1,{_zz_dataShuffle_3_3,_zz_dataShuffle_3_4}}}}}}}}}},_zz_dataShuffle_3[7 : 0]};
      end
      3'b001 : begin
        dataShuffle_3 = {{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_2,{_zz_dataShuffle_3_5,_zz_dataShuffle_3_6}}}}}}}}}},_zz_dataShuffle_3[15 : 0]};
      end
      3'b010 : begin
        dataShuffle_3 = _zz_dataShuffle_3;
      end
      default : begin
        dataShuffle_3 = _zz_dataShuffle_3;
      end
    endcase
  end

  assign _zz_dataShuffle_3_2 = (_zz_dataShuffle_3[15] && stage2In_payload_lsCtrlBundle_signed);
  assign axiShiftedData = (io_axi_rdata >>> missingEntry_vaddr[5 : 0]);
  assign _zz_axiShuffle = (axiShiftedData[7] && stage2In_payload_lsCtrlBundle_signed);
  always @(*) begin
    case(missingEntry_size)
      3'b000 : begin
        axiShuffle = {{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle,{_zz_axiShuffle_2,_zz_axiShuffle_3}}}}}}}}}},axiShiftedData[7 : 0]};
      end
      3'b001 : begin
        axiShuffle = {{_zz_axiShuffle_1,{_zz_axiShuffle_1,{_zz_axiShuffle_1,{_zz_axiShuffle_1,{_zz_axiShuffle_1,{_zz_axiShuffle_1,{_zz_axiShuffle_1,{_zz_axiShuffle_1,{_zz_axiShuffle_1,{_zz_axiShuffle_4,_zz_axiShuffle_5}}}}}}}}}},axiShiftedData[15 : 0]};
      end
      3'b010 : begin
        axiShuffle = axiShiftedData;
      end
      default : begin
        axiShuffle = axiShiftedData;
      end
    endcase
  end

  assign _zz_axiShuffle_1 = (axiShiftedData[15] && stage2In_payload_lsCtrlBundle_signed);
  assign io_output_payload_robIdx = (axiLoad ? missingEntry_robIdx : stage2In_payload_robIdx);
  assign io_output_payload_data = (axiLoad ? (missingEntry_sc ? scResAXI : axiShuffle) : (stage2In_payload_lsCtrlBundle_sc ? scResHit : _zz_io_output_payload_data_3));
  assign io_output_payload_prd = (axiLoad ? missingEntry_prd : stage2In_payload_prd);
  assign io_output_payload_branchResult_targetPC = (axiLoad ? missingEntry_branchResult_targetPC : stage2In_payload_branchResult_targetPC);
  assign io_output_payload_branchResult_branchResult = (axiLoad ? missingEntry_branchResult_branchResult : stage2In_payload_branchResult_branchResult);
  assign io_output_payload_branchResult_predictFail = (axiLoad ? missingEntry_branchResult_predictFail : stage2In_payload_branchResult_predictFail);
  assign io_output_payload_exceptionInfo_exception = (axiLoad ? missingEntry_exceptionInfo_exception : exceptionInfo_exception);
  assign io_output_payload_exceptionInfo_eCode = (axiLoad ? missingEntry_exceptionInfo_eCode : exceptionInfo_eCode);
  assign io_output_payload_exceptionInfo_eSubCode = (axiLoad ? missingEntry_exceptionInfo_eSubCode : exceptionInfo_eSubCode);
  assign io_output_valid = (axiLoad || (((((|hit) || exceptionInfo_exception) || (! stage2In_payload_lsCtrlBundle_normalMemOp)) && stage2In_valid) && (! cacopActive)));
  assign io_badv_robIdx = stage2In_payload_robIdx;
  assign io_badv_vaddr = stage2In_payload_vaddr;
  assign io_badv_wen = (((exceptionInfo_exception && stage2In_valid) && (! cacopActive)) && stage2In_payload_lsException);
  assign io_wakeOut_0_valid = 1'b0;
  assign io_wakeOut_0_payload = 6'h00;
  assign io_wakeOut_1_valid = ((axiCtrl_stateReg == axiCtrl_enumDef_readFirst) || ((((stage2In_valid && (! axiLoad)) && (stage2In_payload_lsCtrlBundle_load || stage2In_payload_lsCtrlBundle_sc)) && (|hit)) && (! cacopActive)));
  assign io_wakeOut_1_payload = io_output_payload_prd;
  assign io_ctrl_busy = ((refilling || rollingBack) || (cacopActive && stage2In_valid));
  assign cacopSetInvalid = (stage2In_payload_isHitInvalidate || stage2In_payload_isIndexInvalidate);
  assign cacopActive = (cacopSetInvalid || stage2In_payload_isStoreTag);
  always @(*) begin
    cacopWriteBack = 1'b0;
    if(when_LSU_l661) begin
      cacopWriteBack = (|wayDirty);
    end
  end

  assign cacopIdx = stage2In_payload_vaddr[10 : 6];
  assign cacopWay = (stage2In_payload_isHitInvalidate ? hit : _zz_cacopWay);
  assign when_LSU_l661 = (stage2In_valid && cacopSetInvalid);
  assign when_LSU_l663 = cacopWay[0];
  assign _zz_61 = ({31'd0,1'b1} <<< cacopIdx);
  assign when_LSU_l663_1 = cacopWay[1];
  assign _zz_62 = ({31'd0,1'b1} <<< cacopIdx);
  assign when_LSU_l663_2 = cacopWay[2];
  assign _zz_63 = ({31'd0,1'b1} <<< cacopIdx);
  assign when_LSU_l663_3 = cacopWay[3];
  assign _zz_64 = ({31'd0,1'b1} <<< cacopIdx);
  assign specialOpBufferWrite = ((((! stage1Out_payload_lsCtrlBundle_normalMemOp) && (io_input_payload_uop_lsuOp != LSUOp_preld)) && (io_input_payload_uop_lsuOp != LSUOp_dbar)) && (! io_ctrl_stall));
  assign io_specialOpBufferUpdate_valid = (io_input_valid && specialOpBufferWrite);
  assign io_specialOpBufferUpdate_payload_uop_lsuOp = io_input_payload_uop_lsuOp;
  assign io_specialOpBufferUpdate_payload_uop_lsuCoOp = io_input_payload_uop_lsuCoOp;
  assign io_specialOpBufferUpdate_payload_vaddr = ((io_input_payload_uop_lsuOp == LSUOp_invtlb) ? io_input_payload_src2 : address);
  assign io_specialOpBufferUpdate_payload_asid = io_input_payload_src1[9 : 0];
  assign io_storeData = stage2In_payload_storeData;
  assign io_storeMask = (stage2In_payload_lsCtrlBundle_store ? stage2In_payload_lsCtrlBundle_lsMask : 4'b0000);
  assign io_VAddr = stage2In_payload_vaddr;
  assign io_PAddr = {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_vaddr[11 : 0]};
  assign io_loadMask = (stage2In_payload_lsCtrlBundle_load ? stage2In_payload_lsCtrlBundle_lsMask : 4'b0000);
  always @(*) begin
    axiCtrl_stateNext = axiCtrl_stateReg;
    case(axiCtrl_stateReg)
      axiCtrl_enumDef_idle : begin
        if(when_LSU_l436) begin
          if(when_LSU_l447) begin
            axiCtrl_stateNext = axiCtrl_enumDef_writeReq;
          end else begin
            axiCtrl_stateNext = axiCtrl_enumDef_readReq;
          end
        end
        if(when_LSU_l453) begin
          axiCtrl_stateNext = axiCtrl_enumDef_writeReq;
        end
      end
      axiCtrl_enumDef_readReq : begin
        if(when_LSU_l480) begin
          if(when_LSU_l481) begin
            axiCtrl_stateNext = axiCtrl_enumDef_readFirst;
          end else begin
            axiCtrl_stateNext = axiCtrl_enumDef_read;
          end
        end
      end
      axiCtrl_enumDef_readFirst : begin
        if(when_LSU_l496) begin
          axiCtrl_stateNext = axiCtrl_enumDef_read;
        end
      end
      axiCtrl_enumDef_read : begin
        if(when_LSU_l510) begin
          if(io_axi_rlast) begin
            axiCtrl_stateNext = axiCtrl_enumDef_idle;
          end
        end
      end
      axiCtrl_enumDef_writeReq : begin
        if(when_LSU_l527) begin
          axiCtrl_stateNext = axiCtrl_enumDef_write;
        end
      end
      axiCtrl_enumDef_write : begin
        if(when_LSU_l539) begin
          if(io_axi_wlast) begin
            if(transferUncached) begin
              axiCtrl_stateNext = axiCtrl_enumDef_idle;
            end else begin
              if(transferCACOP) begin
                axiCtrl_stateNext = axiCtrl_enumDef_idle;
              end else begin
                axiCtrl_stateNext = axiCtrl_enumDef_readReq;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(axiCtrl_wantStart) begin
      axiCtrl_stateNext = axiCtrl_enumDef_idle;
    end
    if(axiCtrl_wantKill) begin
      axiCtrl_stateNext = axiCtrl_enumDef_BOOT;
    end
  end

  assign when_LSU_l436 = ((! io_flush) && (missBufferAllowMask[0] || (missBufferPreAllowMask[0] && (! missingEntry_uncached))));
  assign when_LSU_l447 = ((missingEntry_uncached && missingEntry_store) || missingEntry_writeBack);
  assign when_LSU_l453 = ((cacopSetInvalid && cacopWriteBack) && stage2In_valid);
  assign when_LSU_l471 = (! transferUncached);
  assign when_LSU_l473 = transferWaySelect[0];
  assign _zz_65 = ({31'd0,1'b1} <<< _zz__zz_65[10 : 6]);
  assign _zz_66 = ({31'd0,1'b1} <<< _zz__zz_66[10 : 6]);
  assign when_LSU_l473_1 = transferWaySelect[1];
  assign _zz_67 = ({31'd0,1'b1} <<< _zz__zz_67[10 : 6]);
  assign _zz_68 = ({31'd0,1'b1} <<< _zz__zz_68[10 : 6]);
  assign when_LSU_l473_2 = transferWaySelect[2];
  assign _zz_69 = ({31'd0,1'b1} <<< _zz__zz_69[10 : 6]);
  assign _zz_70 = ({31'd0,1'b1} <<< _zz__zz_70[10 : 6]);
  assign when_LSU_l473_3 = transferWaySelect[3];
  assign _zz_71 = ({31'd0,1'b1} <<< _zz__zz_71[10 : 6]);
  assign _zz_72 = ({31'd0,1'b1} <<< _zz__zz_72[10 : 6]);
  assign when_LSU_l480 = (io_axi_arvalid && io_axi_arready);
  assign when_LSU_l481 = (missingEntry_valid && (! io_flush));
  assign when_LSU_l496 = (io_axi_rvalid && io_axi_rready);
  assign when_LSU_l510 = (io_axi_rvalid && io_axi_rready);
  assign when_LSU_l527 = (io_axi_awvalid && io_axi_awready);
  assign when_LSU_l539 = (io_axi_wvalid && io_axi_wready);
  always @(*) begin
    rollbackCtrl_stateNext = rollbackCtrl_stateReg;
    case(rollbackCtrl_stateReg)
      rollbackCtrl_enumDef_idle : begin
        if(when_LSU_l567) begin
          rollbackCtrl_stateNext = rollbackCtrl_enumDef_rollback;
        end
      end
      rollbackCtrl_enumDef_rollback : begin
        if(when_LSU_l575) begin
          rollbackCtrl_stateNext = rollbackCtrl_enumDef_idle;
        end
      end
      default : begin
      end
    endcase
    if(rollbackCtrl_wantStart) begin
      rollbackCtrl_stateNext = rollbackCtrl_enumDef_idle;
    end
    if(rollbackCtrl_wantKill) begin
      rollbackCtrl_stateNext = rollbackCtrl_enumDef_BOOT;
    end
  end

  assign when_LSU_l564 = (writeBufferAppend && (! io_flush));
  assign when_LSU_l567 = (io_flush && _zz_when_LSU_l567);
  assign when_LSU_l575 = (writeBufferHead == writeBufferTail);
  assign data_0_portA_en = (portRen0_0 && 1'b1);
  assign data_0_portB_en = (portRen1_0 && 1'b1);
  assign data_1_portA_en = (portRen0_1 && 1'b1);
  assign data_1_portB_en = (portRen1_1 && 1'b1);
  assign data_2_portA_en = (portRen0_2 && 1'b1);
  assign data_2_portB_en = (portRen1_2 && 1'b1);
  assign data_3_portA_en = (portRen0_3 && 1'b1);
  assign data_3_portB_en = (portRen1_3 && 1'b1);
  assign tag_0_wr_en = (_zz_wr_en_3 && 1'b1);
  assign tag_0_wr_addr = _zz_wr_addr[10 : 6];
  assign tag_0_wr_data = {stage2In_payload_tlb_pageInfo_ppn,_zz_wr_data[11 : 11]};
  assign tag_0_wr_mask = 1'b1;
  assign tag_0_rd_en = (stage1Out_fire && 1'b1);
  assign tag_0_rd_addr = _zz_rd_addr[10 : 6];
  assign tag_1_wr_en = (_zz_wr_en_2 && 1'b1);
  assign tag_1_wr_addr = _zz_wr_addr_1[10 : 6];
  assign tag_1_wr_data = {stage2In_payload_tlb_pageInfo_ppn,_zz_wr_data_1[11 : 11]};
  assign tag_1_wr_mask = 1'b1;
  assign tag_1_rd_en = (stage1Out_fire && 1'b1);
  assign tag_1_rd_addr = _zz_rd_addr_1[10 : 6];
  assign tag_2_wr_en = (_zz_wr_en_1 && 1'b1);
  assign tag_2_wr_addr = _zz_wr_addr_2[10 : 6];
  assign tag_2_wr_data = {stage2In_payload_tlb_pageInfo_ppn,_zz_wr_data_2[11 : 11]};
  assign tag_2_wr_mask = 1'b1;
  assign tag_2_rd_en = (stage1Out_fire && 1'b1);
  assign tag_2_rd_addr = _zz_rd_addr_2[10 : 6];
  assign tag_3_wr_en = (_zz_wr_en && 1'b1);
  assign tag_3_wr_addr = _zz_wr_addr_3[10 : 6];
  assign tag_3_wr_data = {stage2In_payload_tlb_pageInfo_ppn,_zz_wr_data_3[11 : 11]};
  assign tag_3_wr_mask = 1'b1;
  assign tag_3_rd_en = (stage1Out_fire && 1'b1);
  assign tag_3_rd_addr = _zz_rd_addr_3[10 : 6];
  always @(posedge aclk) begin
    if(!aresetn) begin
      valid_0_0 <= 1'b0;
      valid_0_1 <= 1'b0;
      valid_0_2 <= 1'b0;
      valid_0_3 <= 1'b0;
      valid_0_4 <= 1'b0;
      valid_0_5 <= 1'b0;
      valid_0_6 <= 1'b0;
      valid_0_7 <= 1'b0;
      valid_0_8 <= 1'b0;
      valid_0_9 <= 1'b0;
      valid_0_10 <= 1'b0;
      valid_0_11 <= 1'b0;
      valid_0_12 <= 1'b0;
      valid_0_13 <= 1'b0;
      valid_0_14 <= 1'b0;
      valid_0_15 <= 1'b0;
      valid_0_16 <= 1'b0;
      valid_0_17 <= 1'b0;
      valid_0_18 <= 1'b0;
      valid_0_19 <= 1'b0;
      valid_0_20 <= 1'b0;
      valid_0_21 <= 1'b0;
      valid_0_22 <= 1'b0;
      valid_0_23 <= 1'b0;
      valid_0_24 <= 1'b0;
      valid_0_25 <= 1'b0;
      valid_0_26 <= 1'b0;
      valid_0_27 <= 1'b0;
      valid_0_28 <= 1'b0;
      valid_0_29 <= 1'b0;
      valid_0_30 <= 1'b0;
      valid_0_31 <= 1'b0;
      valid_1_0 <= 1'b0;
      valid_1_1 <= 1'b0;
      valid_1_2 <= 1'b0;
      valid_1_3 <= 1'b0;
      valid_1_4 <= 1'b0;
      valid_1_5 <= 1'b0;
      valid_1_6 <= 1'b0;
      valid_1_7 <= 1'b0;
      valid_1_8 <= 1'b0;
      valid_1_9 <= 1'b0;
      valid_1_10 <= 1'b0;
      valid_1_11 <= 1'b0;
      valid_1_12 <= 1'b0;
      valid_1_13 <= 1'b0;
      valid_1_14 <= 1'b0;
      valid_1_15 <= 1'b0;
      valid_1_16 <= 1'b0;
      valid_1_17 <= 1'b0;
      valid_1_18 <= 1'b0;
      valid_1_19 <= 1'b0;
      valid_1_20 <= 1'b0;
      valid_1_21 <= 1'b0;
      valid_1_22 <= 1'b0;
      valid_1_23 <= 1'b0;
      valid_1_24 <= 1'b0;
      valid_1_25 <= 1'b0;
      valid_1_26 <= 1'b0;
      valid_1_27 <= 1'b0;
      valid_1_28 <= 1'b0;
      valid_1_29 <= 1'b0;
      valid_1_30 <= 1'b0;
      valid_1_31 <= 1'b0;
      valid_2_0 <= 1'b0;
      valid_2_1 <= 1'b0;
      valid_2_2 <= 1'b0;
      valid_2_3 <= 1'b0;
      valid_2_4 <= 1'b0;
      valid_2_5 <= 1'b0;
      valid_2_6 <= 1'b0;
      valid_2_7 <= 1'b0;
      valid_2_8 <= 1'b0;
      valid_2_9 <= 1'b0;
      valid_2_10 <= 1'b0;
      valid_2_11 <= 1'b0;
      valid_2_12 <= 1'b0;
      valid_2_13 <= 1'b0;
      valid_2_14 <= 1'b0;
      valid_2_15 <= 1'b0;
      valid_2_16 <= 1'b0;
      valid_2_17 <= 1'b0;
      valid_2_18 <= 1'b0;
      valid_2_19 <= 1'b0;
      valid_2_20 <= 1'b0;
      valid_2_21 <= 1'b0;
      valid_2_22 <= 1'b0;
      valid_2_23 <= 1'b0;
      valid_2_24 <= 1'b0;
      valid_2_25 <= 1'b0;
      valid_2_26 <= 1'b0;
      valid_2_27 <= 1'b0;
      valid_2_28 <= 1'b0;
      valid_2_29 <= 1'b0;
      valid_2_30 <= 1'b0;
      valid_2_31 <= 1'b0;
      valid_3_0 <= 1'b0;
      valid_3_1 <= 1'b0;
      valid_3_2 <= 1'b0;
      valid_3_3 <= 1'b0;
      valid_3_4 <= 1'b0;
      valid_3_5 <= 1'b0;
      valid_3_6 <= 1'b0;
      valid_3_7 <= 1'b0;
      valid_3_8 <= 1'b0;
      valid_3_9 <= 1'b0;
      valid_3_10 <= 1'b0;
      valid_3_11 <= 1'b0;
      valid_3_12 <= 1'b0;
      valid_3_13 <= 1'b0;
      valid_3_14 <= 1'b0;
      valid_3_15 <= 1'b0;
      valid_3_16 <= 1'b0;
      valid_3_17 <= 1'b0;
      valid_3_18 <= 1'b0;
      valid_3_19 <= 1'b0;
      valid_3_20 <= 1'b0;
      valid_3_21 <= 1'b0;
      valid_3_22 <= 1'b0;
      valid_3_23 <= 1'b0;
      valid_3_24 <= 1'b0;
      valid_3_25 <= 1'b0;
      valid_3_26 <= 1'b0;
      valid_3_27 <= 1'b0;
      valid_3_28 <= 1'b0;
      valid_3_29 <= 1'b0;
      valid_3_30 <= 1'b0;
      valid_3_31 <= 1'b0;
      dirty_0_0 <= 1'b0;
      dirty_0_1 <= 1'b0;
      dirty_0_2 <= 1'b0;
      dirty_0_3 <= 1'b0;
      dirty_0_4 <= 1'b0;
      dirty_0_5 <= 1'b0;
      dirty_0_6 <= 1'b0;
      dirty_0_7 <= 1'b0;
      dirty_0_8 <= 1'b0;
      dirty_0_9 <= 1'b0;
      dirty_0_10 <= 1'b0;
      dirty_0_11 <= 1'b0;
      dirty_0_12 <= 1'b0;
      dirty_0_13 <= 1'b0;
      dirty_0_14 <= 1'b0;
      dirty_0_15 <= 1'b0;
      dirty_0_16 <= 1'b0;
      dirty_0_17 <= 1'b0;
      dirty_0_18 <= 1'b0;
      dirty_0_19 <= 1'b0;
      dirty_0_20 <= 1'b0;
      dirty_0_21 <= 1'b0;
      dirty_0_22 <= 1'b0;
      dirty_0_23 <= 1'b0;
      dirty_0_24 <= 1'b0;
      dirty_0_25 <= 1'b0;
      dirty_0_26 <= 1'b0;
      dirty_0_27 <= 1'b0;
      dirty_0_28 <= 1'b0;
      dirty_0_29 <= 1'b0;
      dirty_0_30 <= 1'b0;
      dirty_0_31 <= 1'b0;
      dirty_1_0 <= 1'b0;
      dirty_1_1 <= 1'b0;
      dirty_1_2 <= 1'b0;
      dirty_1_3 <= 1'b0;
      dirty_1_4 <= 1'b0;
      dirty_1_5 <= 1'b0;
      dirty_1_6 <= 1'b0;
      dirty_1_7 <= 1'b0;
      dirty_1_8 <= 1'b0;
      dirty_1_9 <= 1'b0;
      dirty_1_10 <= 1'b0;
      dirty_1_11 <= 1'b0;
      dirty_1_12 <= 1'b0;
      dirty_1_13 <= 1'b0;
      dirty_1_14 <= 1'b0;
      dirty_1_15 <= 1'b0;
      dirty_1_16 <= 1'b0;
      dirty_1_17 <= 1'b0;
      dirty_1_18 <= 1'b0;
      dirty_1_19 <= 1'b0;
      dirty_1_20 <= 1'b0;
      dirty_1_21 <= 1'b0;
      dirty_1_22 <= 1'b0;
      dirty_1_23 <= 1'b0;
      dirty_1_24 <= 1'b0;
      dirty_1_25 <= 1'b0;
      dirty_1_26 <= 1'b0;
      dirty_1_27 <= 1'b0;
      dirty_1_28 <= 1'b0;
      dirty_1_29 <= 1'b0;
      dirty_1_30 <= 1'b0;
      dirty_1_31 <= 1'b0;
      dirty_2_0 <= 1'b0;
      dirty_2_1 <= 1'b0;
      dirty_2_2 <= 1'b0;
      dirty_2_3 <= 1'b0;
      dirty_2_4 <= 1'b0;
      dirty_2_5 <= 1'b0;
      dirty_2_6 <= 1'b0;
      dirty_2_7 <= 1'b0;
      dirty_2_8 <= 1'b0;
      dirty_2_9 <= 1'b0;
      dirty_2_10 <= 1'b0;
      dirty_2_11 <= 1'b0;
      dirty_2_12 <= 1'b0;
      dirty_2_13 <= 1'b0;
      dirty_2_14 <= 1'b0;
      dirty_2_15 <= 1'b0;
      dirty_2_16 <= 1'b0;
      dirty_2_17 <= 1'b0;
      dirty_2_18 <= 1'b0;
      dirty_2_19 <= 1'b0;
      dirty_2_20 <= 1'b0;
      dirty_2_21 <= 1'b0;
      dirty_2_22 <= 1'b0;
      dirty_2_23 <= 1'b0;
      dirty_2_24 <= 1'b0;
      dirty_2_25 <= 1'b0;
      dirty_2_26 <= 1'b0;
      dirty_2_27 <= 1'b0;
      dirty_2_28 <= 1'b0;
      dirty_2_29 <= 1'b0;
      dirty_2_30 <= 1'b0;
      dirty_2_31 <= 1'b0;
      dirty_3_0 <= 1'b0;
      dirty_3_1 <= 1'b0;
      dirty_3_2 <= 1'b0;
      dirty_3_3 <= 1'b0;
      dirty_3_4 <= 1'b0;
      dirty_3_5 <= 1'b0;
      dirty_3_6 <= 1'b0;
      dirty_3_7 <= 1'b0;
      dirty_3_8 <= 1'b0;
      dirty_3_9 <= 1'b0;
      dirty_3_10 <= 1'b0;
      dirty_3_11 <= 1'b0;
      dirty_3_12 <= 1'b0;
      dirty_3_13 <= 1'b0;
      dirty_3_14 <= 1'b0;
      dirty_3_15 <= 1'b0;
      dirty_3_16 <= 1'b0;
      dirty_3_17 <= 1'b0;
      dirty_3_18 <= 1'b0;
      dirty_3_19 <= 1'b0;
      dirty_3_20 <= 1'b0;
      dirty_3_21 <= 1'b0;
      dirty_3_22 <= 1'b0;
      dirty_3_23 <= 1'b0;
      dirty_3_24 <= 1'b0;
      dirty_3_25 <= 1'b0;
      dirty_3_26 <= 1'b0;
      dirty_3_27 <= 1'b0;
      dirty_3_28 <= 1'b0;
      dirty_3_29 <= 1'b0;
      dirty_3_30 <= 1'b0;
      dirty_3_31 <= 1'b0;
      wayDirtyBypass <= 4'b0000;
      stage1Out_thrown_rValid <= 1'b0;
      transferRAddrHi <= 26'h0000000;
      transferRAddrMid <= 4'b0000;
      transferRAddrLo <= 2'b00;
      transferWAddrHi <= 26'h0000000;
      transferWAddrMid <= 4'b0000;
      transferWAddrLo <= 2'b00;
      transferUncached <= 1'b0;
      transferCACOP <= 1'b0;
      transferWData <= 32'h00000000;
      transferLSMask <= 4'b0000;
      transferWaySelect <= 4'b0000;
      portWData1Bypass_0 <= 32'h00000000;
      portWMask1Bypass_0 <= 4'b0000;
      portWData1Bypass_1 <= 32'h00000000;
      portWMask1Bypass_1 <= 4'b0000;
      portWData1Bypass_2 <= 32'h00000000;
      portWMask1Bypass_2 <= 4'b0000;
      portWData1Bypass_3 <= 32'h00000000;
      portWMask1Bypass_3 <= 4'b0000;
      writeBufferHead <= 3'b000;
      writeBufferTail <= 3'b000;
      writeBuffer_0_robIdx <= 5'h00;
      writeBuffer_0_waySelect <= 4'b0000;
      writeBuffer_0_prevData <= 32'h00000000;
      writeBuffer_0_prevDirty <= 1'b0;
      writeBuffer_0_index <= 9'h000;
      writeBuffer_0_miss <= 1'b0;
      writeBuffer_0_valid <= 1'b0;
      writeBuffer_1_robIdx <= 5'h00;
      writeBuffer_1_waySelect <= 4'b0000;
      writeBuffer_1_prevData <= 32'h00000000;
      writeBuffer_1_prevDirty <= 1'b0;
      writeBuffer_1_index <= 9'h000;
      writeBuffer_1_miss <= 1'b0;
      writeBuffer_1_valid <= 1'b0;
      writeBuffer_2_robIdx <= 5'h00;
      writeBuffer_2_waySelect <= 4'b0000;
      writeBuffer_2_prevData <= 32'h00000000;
      writeBuffer_2_prevDirty <= 1'b0;
      writeBuffer_2_index <= 9'h000;
      writeBuffer_2_miss <= 1'b0;
      writeBuffer_2_valid <= 1'b0;
      writeBuffer_3_robIdx <= 5'h00;
      writeBuffer_3_waySelect <= 4'b0000;
      writeBuffer_3_prevData <= 32'h00000000;
      writeBuffer_3_prevDirty <= 1'b0;
      writeBuffer_3_index <= 9'h000;
      writeBuffer_3_miss <= 1'b0;
      writeBuffer_3_valid <= 1'b0;
      writeBuffer_4_robIdx <= 5'h00;
      writeBuffer_4_waySelect <= 4'b0000;
      writeBuffer_4_prevData <= 32'h00000000;
      writeBuffer_4_prevDirty <= 1'b0;
      writeBuffer_4_index <= 9'h000;
      writeBuffer_4_miss <= 1'b0;
      writeBuffer_4_valid <= 1'b0;
      writeBuffer_5_robIdx <= 5'h00;
      writeBuffer_5_waySelect <= 4'b0000;
      writeBuffer_5_prevData <= 32'h00000000;
      writeBuffer_5_prevDirty <= 1'b0;
      writeBuffer_5_index <= 9'h000;
      writeBuffer_5_miss <= 1'b0;
      writeBuffer_5_valid <= 1'b0;
      writeBuffer_6_robIdx <= 5'h00;
      writeBuffer_6_waySelect <= 4'b0000;
      writeBuffer_6_prevData <= 32'h00000000;
      writeBuffer_6_prevDirty <= 1'b0;
      writeBuffer_6_index <= 9'h000;
      writeBuffer_6_miss <= 1'b0;
      writeBuffer_6_valid <= 1'b0;
      writeBuffer_7_robIdx <= 5'h00;
      writeBuffer_7_waySelect <= 4'b0000;
      writeBuffer_7_prevData <= 32'h00000000;
      writeBuffer_7_prevDirty <= 1'b0;
      writeBuffer_7_index <= 9'h000;
      writeBuffer_7_miss <= 1'b0;
      writeBuffer_7_valid <= 1'b0;
      missBuffer_0_robIdx <= 5'h00;
      missBuffer_0_prd <= 6'h00;
      missBuffer_0_branchResult_targetPC <= 32'h00000000;
      missBuffer_0_branchResult_branchResult <= 1'b0;
      missBuffer_0_branchResult_predictFail <= 1'b0;
      missBuffer_0_exceptionInfo_exception <= 1'b0;
      missBuffer_0_exceptionInfo_eCode <= 6'h00;
      missBuffer_0_exceptionInfo_eSubCode <= 1'b0;
      missBuffer_0_uncached <= 1'b0;
      missBuffer_0_load <= 1'b0;
      missBuffer_0_store <= 1'b0;
      missBuffer_0_signed <= 1'b0;
      missBuffer_0_ll <= 1'b0;
      missBuffer_0_sc <= 1'b0;
      missBuffer_0_writeBufferIdx <= 3'b000;
      missBuffer_0_waySelect <= 4'b0000;
      missBuffer_0_writeBack <= 1'b0;
      missBuffer_0_storeData <= 32'h00000000;
      missBuffer_0_lsMask <= 4'b0000;
      missBuffer_0_size <= 3'b000;
      missBuffer_0_vaddr <= 32'h00000000;
      missBuffer_0_paddr <= 32'h00000000;
      missBuffer_0_prevPaddr <= 32'h00000000;
      missBuffer_0_valid <= 1'b0;
      lruBit_0_0 <= 1'b0;
      lruBit_0_1 <= 1'b0;
      lruBit_0_2 <= 1'b0;
      lruBit_1_0 <= 1'b0;
      lruBit_1_1 <= 1'b0;
      lruBit_1_2 <= 1'b0;
      lruBit_2_0 <= 1'b0;
      lruBit_2_1 <= 1'b0;
      lruBit_2_2 <= 1'b0;
      lruBit_3_0 <= 1'b0;
      lruBit_3_1 <= 1'b0;
      lruBit_3_2 <= 1'b0;
      lruBit_4_0 <= 1'b0;
      lruBit_4_1 <= 1'b0;
      lruBit_4_2 <= 1'b0;
      lruBit_5_0 <= 1'b0;
      lruBit_5_1 <= 1'b0;
      lruBit_5_2 <= 1'b0;
      lruBit_6_0 <= 1'b0;
      lruBit_6_1 <= 1'b0;
      lruBit_6_2 <= 1'b0;
      lruBit_7_0 <= 1'b0;
      lruBit_7_1 <= 1'b0;
      lruBit_7_2 <= 1'b0;
      lruBit_8_0 <= 1'b0;
      lruBit_8_1 <= 1'b0;
      lruBit_8_2 <= 1'b0;
      lruBit_9_0 <= 1'b0;
      lruBit_9_1 <= 1'b0;
      lruBit_9_2 <= 1'b0;
      lruBit_10_0 <= 1'b0;
      lruBit_10_1 <= 1'b0;
      lruBit_10_2 <= 1'b0;
      lruBit_11_0 <= 1'b0;
      lruBit_11_1 <= 1'b0;
      lruBit_11_2 <= 1'b0;
      lruBit_12_0 <= 1'b0;
      lruBit_12_1 <= 1'b0;
      lruBit_12_2 <= 1'b0;
      lruBit_13_0 <= 1'b0;
      lruBit_13_1 <= 1'b0;
      lruBit_13_2 <= 1'b0;
      lruBit_14_0 <= 1'b0;
      lruBit_14_1 <= 1'b0;
      lruBit_14_2 <= 1'b0;
      lruBit_15_0 <= 1'b0;
      lruBit_15_1 <= 1'b0;
      lruBit_15_2 <= 1'b0;
      lruBit_16_0 <= 1'b0;
      lruBit_16_1 <= 1'b0;
      lruBit_16_2 <= 1'b0;
      lruBit_17_0 <= 1'b0;
      lruBit_17_1 <= 1'b0;
      lruBit_17_2 <= 1'b0;
      lruBit_18_0 <= 1'b0;
      lruBit_18_1 <= 1'b0;
      lruBit_18_2 <= 1'b0;
      lruBit_19_0 <= 1'b0;
      lruBit_19_1 <= 1'b0;
      lruBit_19_2 <= 1'b0;
      lruBit_20_0 <= 1'b0;
      lruBit_20_1 <= 1'b0;
      lruBit_20_2 <= 1'b0;
      lruBit_21_0 <= 1'b0;
      lruBit_21_1 <= 1'b0;
      lruBit_21_2 <= 1'b0;
      lruBit_22_0 <= 1'b0;
      lruBit_22_1 <= 1'b0;
      lruBit_22_2 <= 1'b0;
      lruBit_23_0 <= 1'b0;
      lruBit_23_1 <= 1'b0;
      lruBit_23_2 <= 1'b0;
      lruBit_24_0 <= 1'b0;
      lruBit_24_1 <= 1'b0;
      lruBit_24_2 <= 1'b0;
      lruBit_25_0 <= 1'b0;
      lruBit_25_1 <= 1'b0;
      lruBit_25_2 <= 1'b0;
      lruBit_26_0 <= 1'b0;
      lruBit_26_1 <= 1'b0;
      lruBit_26_2 <= 1'b0;
      lruBit_27_0 <= 1'b0;
      lruBit_27_1 <= 1'b0;
      lruBit_27_2 <= 1'b0;
      lruBit_28_0 <= 1'b0;
      lruBit_28_1 <= 1'b0;
      lruBit_28_2 <= 1'b0;
      lruBit_29_0 <= 1'b0;
      lruBit_29_1 <= 1'b0;
      lruBit_29_2 <= 1'b0;
      lruBit_30_0 <= 1'b0;
      lruBit_30_1 <= 1'b0;
      lruBit_30_2 <= 1'b0;
      lruBit_31_0 <= 1'b0;
      lruBit_31_1 <= 1'b0;
      lruBit_31_2 <= 1'b0;
      axiCtrl_stateReg <= axiCtrl_enumDef_BOOT;
      rollbackCtrl_stateReg <= rollbackCtrl_enumDef_BOOT;
    end else begin
      if(stage1Out_thrown_ready) begin
        stage1Out_thrown_rValid <= stage1Out_thrown_valid;
      end
      if(portRen0_0) begin
        if(when_LSU_l174) begin
          portWData1Bypass_0 <= portWData1;
          portWMask1Bypass_0 <= portWMask1;
        end else begin
          portWData1Bypass_0 <= 32'h00000000;
          portWMask1Bypass_0 <= 4'b0000;
        end
      end
      if(portRen0_1) begin
        if(when_LSU_l174_1) begin
          portWData1Bypass_1 <= portWData1;
          portWMask1Bypass_1 <= portWMask1;
        end else begin
          portWData1Bypass_1 <= 32'h00000000;
          portWMask1Bypass_1 <= 4'b0000;
        end
      end
      if(portRen0_2) begin
        if(when_LSU_l174_2) begin
          portWData1Bypass_2 <= portWData1;
          portWMask1Bypass_2 <= portWMask1;
        end else begin
          portWData1Bypass_2 <= 32'h00000000;
          portWMask1Bypass_2 <= 4'b0000;
        end
      end
      if(portRen0_3) begin
        if(when_LSU_l174_3) begin
          portWData1Bypass_3 <= portWData1;
          portWMask1Bypass_3 <= portWMask1;
        end else begin
          portWData1Bypass_3 <= 32'h00000000;
          portWMask1Bypass_3 <= 4'b0000;
        end
      end
      writeBufferHead <= writeBufferHeadNext;
      if(when_LSU_l267) begin
        if(_zz_2) begin
          writeBuffer_0_robIdx <= stage2In_payload_robIdx;
        end
        if(_zz_3) begin
          writeBuffer_1_robIdx <= stage2In_payload_robIdx;
        end
        if(_zz_4) begin
          writeBuffer_2_robIdx <= stage2In_payload_robIdx;
        end
        if(_zz_5) begin
          writeBuffer_3_robIdx <= stage2In_payload_robIdx;
        end
        if(_zz_6) begin
          writeBuffer_4_robIdx <= stage2In_payload_robIdx;
        end
        if(_zz_7) begin
          writeBuffer_5_robIdx <= stage2In_payload_robIdx;
        end
        if(_zz_8) begin
          writeBuffer_6_robIdx <= stage2In_payload_robIdx;
        end
        if(_zz_9) begin
          writeBuffer_7_robIdx <= stage2In_payload_robIdx;
        end
        if(_zz_2) begin
          writeBuffer_0_waySelect <= _zz_writeBuffer_0_waySelect;
        end
        if(_zz_3) begin
          writeBuffer_1_waySelect <= _zz_writeBuffer_0_waySelect;
        end
        if(_zz_4) begin
          writeBuffer_2_waySelect <= _zz_writeBuffer_0_waySelect;
        end
        if(_zz_5) begin
          writeBuffer_3_waySelect <= _zz_writeBuffer_0_waySelect;
        end
        if(_zz_6) begin
          writeBuffer_4_waySelect <= _zz_writeBuffer_0_waySelect;
        end
        if(_zz_7) begin
          writeBuffer_5_waySelect <= _zz_writeBuffer_0_waySelect;
        end
        if(_zz_8) begin
          writeBuffer_6_waySelect <= _zz_writeBuffer_0_waySelect;
        end
        if(_zz_9) begin
          writeBuffer_7_waySelect <= _zz_writeBuffer_0_waySelect;
        end
        if(_zz_2) begin
          writeBuffer_0_prevData <= _zz_writeBuffer_0_prevData;
        end
        if(_zz_3) begin
          writeBuffer_1_prevData <= _zz_writeBuffer_0_prevData;
        end
        if(_zz_4) begin
          writeBuffer_2_prevData <= _zz_writeBuffer_0_prevData;
        end
        if(_zz_5) begin
          writeBuffer_3_prevData <= _zz_writeBuffer_0_prevData;
        end
        if(_zz_6) begin
          writeBuffer_4_prevData <= _zz_writeBuffer_0_prevData;
        end
        if(_zz_7) begin
          writeBuffer_5_prevData <= _zz_writeBuffer_0_prevData;
        end
        if(_zz_8) begin
          writeBuffer_6_prevData <= _zz_writeBuffer_0_prevData;
        end
        if(_zz_9) begin
          writeBuffer_7_prevData <= _zz_writeBuffer_0_prevData;
        end
        if(_zz_2) begin
          writeBuffer_0_prevDirty <= _zz_writeBuffer_0_prevDirty;
        end
        if(_zz_3) begin
          writeBuffer_1_prevDirty <= _zz_writeBuffer_0_prevDirty;
        end
        if(_zz_4) begin
          writeBuffer_2_prevDirty <= _zz_writeBuffer_0_prevDirty;
        end
        if(_zz_5) begin
          writeBuffer_3_prevDirty <= _zz_writeBuffer_0_prevDirty;
        end
        if(_zz_6) begin
          writeBuffer_4_prevDirty <= _zz_writeBuffer_0_prevDirty;
        end
        if(_zz_7) begin
          writeBuffer_5_prevDirty <= _zz_writeBuffer_0_prevDirty;
        end
        if(_zz_8) begin
          writeBuffer_6_prevDirty <= _zz_writeBuffer_0_prevDirty;
        end
        if(_zz_9) begin
          writeBuffer_7_prevDirty <= _zz_writeBuffer_0_prevDirty;
        end
        if(_zz_2) begin
          writeBuffer_0_index <= _zz_writeBuffer_0_index;
        end
        if(_zz_3) begin
          writeBuffer_1_index <= _zz_writeBuffer_0_index;
        end
        if(_zz_4) begin
          writeBuffer_2_index <= _zz_writeBuffer_0_index;
        end
        if(_zz_5) begin
          writeBuffer_3_index <= _zz_writeBuffer_0_index;
        end
        if(_zz_6) begin
          writeBuffer_4_index <= _zz_writeBuffer_0_index;
        end
        if(_zz_7) begin
          writeBuffer_5_index <= _zz_writeBuffer_0_index;
        end
        if(_zz_8) begin
          writeBuffer_6_index <= _zz_writeBuffer_0_index;
        end
        if(_zz_9) begin
          writeBuffer_7_index <= _zz_writeBuffer_0_index;
        end
        if(_zz_2) begin
          writeBuffer_0_miss <= miss;
        end
        if(_zz_3) begin
          writeBuffer_1_miss <= miss;
        end
        if(_zz_4) begin
          writeBuffer_2_miss <= miss;
        end
        if(_zz_5) begin
          writeBuffer_3_miss <= miss;
        end
        if(_zz_6) begin
          writeBuffer_4_miss <= miss;
        end
        if(_zz_7) begin
          writeBuffer_5_miss <= miss;
        end
        if(_zz_8) begin
          writeBuffer_6_miss <= miss;
        end
        if(_zz_9) begin
          writeBuffer_7_miss <= miss;
        end
      end
      if(writeBufferUpdate) begin
        if(_zz_11) begin
          writeBuffer_0_prevData <= io_axi_rdata;
        end
        if(_zz_12) begin
          writeBuffer_1_prevData <= io_axi_rdata;
        end
        if(_zz_13) begin
          writeBuffer_2_prevData <= io_axi_rdata;
        end
        if(_zz_14) begin
          writeBuffer_3_prevData <= io_axi_rdata;
        end
        if(_zz_15) begin
          writeBuffer_4_prevData <= io_axi_rdata;
        end
        if(_zz_16) begin
          writeBuffer_5_prevData <= io_axi_rdata;
        end
        if(_zz_17) begin
          writeBuffer_6_prevData <= io_axi_rdata;
        end
        if(_zz_18) begin
          writeBuffer_7_prevData <= io_axi_rdata;
        end
        if(_zz_11) begin
          writeBuffer_0_miss <= 1'b0;
        end
        if(_zz_12) begin
          writeBuffer_1_miss <= 1'b0;
        end
        if(_zz_13) begin
          writeBuffer_2_miss <= 1'b0;
        end
        if(_zz_14) begin
          writeBuffer_3_miss <= 1'b0;
        end
        if(_zz_15) begin
          writeBuffer_4_miss <= 1'b0;
        end
        if(_zz_16) begin
          writeBuffer_5_miss <= 1'b0;
        end
        if(_zz_17) begin
          writeBuffer_6_miss <= 1'b0;
        end
        if(_zz_18) begin
          writeBuffer_7_miss <= 1'b0;
        end
      end
      writeBuffer_0_valid <= ((writeBufferRetireMask[0] || (rollingBack && (writeBufferTail == 3'b000))) ? 1'b0 : (writeBuffer_0_valid || ((writeBufferAppend && (writeBufferTail == 3'b000)) && (! io_flush))));
      writeBuffer_1_valid <= ((writeBufferRetireMask[1] || (rollingBack && (writeBufferTail == 3'b001))) ? 1'b0 : (writeBuffer_1_valid || ((writeBufferAppend && (writeBufferTail == 3'b001)) && (! io_flush))));
      writeBuffer_2_valid <= ((writeBufferRetireMask[2] || (rollingBack && (writeBufferTail == 3'b010))) ? 1'b0 : (writeBuffer_2_valid || ((writeBufferAppend && (writeBufferTail == 3'b010)) && (! io_flush))));
      writeBuffer_3_valid <= ((writeBufferRetireMask[3] || (rollingBack && (writeBufferTail == 3'b011))) ? 1'b0 : (writeBuffer_3_valid || ((writeBufferAppend && (writeBufferTail == 3'b011)) && (! io_flush))));
      writeBuffer_4_valid <= ((writeBufferRetireMask[4] || (rollingBack && (writeBufferTail == 3'b100))) ? 1'b0 : (writeBuffer_4_valid || ((writeBufferAppend && (writeBufferTail == 3'b100)) && (! io_flush))));
      writeBuffer_5_valid <= ((writeBufferRetireMask[5] || (rollingBack && (writeBufferTail == 3'b101))) ? 1'b0 : (writeBuffer_5_valid || ((writeBufferAppend && (writeBufferTail == 3'b101)) && (! io_flush))));
      writeBuffer_6_valid <= ((writeBufferRetireMask[6] || (rollingBack && (writeBufferTail == 3'b110))) ? 1'b0 : (writeBuffer_6_valid || ((writeBufferAppend && (writeBufferTail == 3'b110)) && (! io_flush))));
      writeBuffer_7_valid <= ((writeBufferRetireMask[7] || (rollingBack && (writeBufferTail == 3'b111))) ? 1'b0 : (writeBuffer_7_valid || ((writeBufferAppend && (writeBufferTail == 3'b111)) && (! io_flush))));
      if(when_LSU_l292) begin
        if(_zz_19) begin
          missBuffer_0_robIdx <= stage2In_payload_robIdx;
        end
        if(_zz_19) begin
          missBuffer_0_prd <= stage2In_payload_prd;
        end
        if(_zz_19) begin
          missBuffer_0_branchResult_targetPC <= stage2In_payload_branchResult_targetPC;
        end
        if(_zz_19) begin
          missBuffer_0_branchResult_branchResult <= stage2In_payload_branchResult_branchResult;
        end
        if(_zz_19) begin
          missBuffer_0_branchResult_predictFail <= stage2In_payload_branchResult_predictFail;
        end
        if(_zz_19) begin
          missBuffer_0_exceptionInfo_exception <= exceptionInfo_exception;
        end
        if(_zz_19) begin
          missBuffer_0_exceptionInfo_eCode <= exceptionInfo_eCode;
        end
        if(_zz_19) begin
          missBuffer_0_exceptionInfo_eSubCode <= exceptionInfo_eSubCode;
        end
        if(_zz_19) begin
          missBuffer_0_uncached <= (stage2In_payload_tlb_pageInfo_mat == 2'b00);
        end
        if(_zz_19) begin
          missBuffer_0_load <= stage2In_payload_lsCtrlBundle_load;
        end
        if(_zz_19) begin
          missBuffer_0_store <= stage2In_payload_lsCtrlBundle_store;
        end
        if(_zz_19) begin
          missBuffer_0_signed <= stage2In_payload_lsCtrlBundle_signed;
        end
        if(_zz_19) begin
          missBuffer_0_ll <= stage2In_payload_lsCtrlBundle_ll;
        end
        if(_zz_19) begin
          missBuffer_0_sc <= stage2In_payload_lsCtrlBundle_sc;
        end
        if(_zz_19) begin
          missBuffer_0_writeBufferIdx <= writeBufferTail;
        end
        if(_zz_19) begin
          missBuffer_0_waySelect <= wayToReplace;
        end
        if(_zz_19) begin
          missBuffer_0_writeBack <= _zz_missBuffer_0_writeBack_8;
        end
        if(_zz_19) begin
          missBuffer_0_storeData <= stage2In_payload_storeData;
        end
        if(_zz_19) begin
          missBuffer_0_lsMask <= realLSMask;
        end
        if(_zz_19) begin
          missBuffer_0_size <= stage2In_payload_lsCtrlBundle_size;
        end
        if(_zz_19) begin
          missBuffer_0_vaddr <= stage2In_payload_vaddr;
        end
        if(_zz_19) begin
          missBuffer_0_paddr <= {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_vaddr[11 : 0]};
        end
        if(_zz_19) begin
          missBuffer_0_prevPaddr <= {_zz_missBuffer_0_prevPaddr,stage2In_payload_vaddr[10 : 0]};
        end
      end
      missBuffer_0_valid <= ((io_flush || (axiFinish && 1'b1)) ? 1'b0 : (missBuffer_0_valid || ((miss && stage2In_ready) && 1'b1)));
      if(when_LSU_l335) begin
        if(_zz_21) begin
          lruBit_0_0 <= _zz_lruBit_0_0;
        end
        if(_zz_22) begin
          lruBit_1_0 <= _zz_lruBit_0_0;
        end
        if(_zz_23) begin
          lruBit_2_0 <= _zz_lruBit_0_0;
        end
        if(_zz_24) begin
          lruBit_3_0 <= _zz_lruBit_0_0;
        end
        if(_zz_25) begin
          lruBit_4_0 <= _zz_lruBit_0_0;
        end
        if(_zz_26) begin
          lruBit_5_0 <= _zz_lruBit_0_0;
        end
        if(_zz_27) begin
          lruBit_6_0 <= _zz_lruBit_0_0;
        end
        if(_zz_28) begin
          lruBit_7_0 <= _zz_lruBit_0_0;
        end
        if(_zz_29) begin
          lruBit_8_0 <= _zz_lruBit_0_0;
        end
        if(_zz_30) begin
          lruBit_9_0 <= _zz_lruBit_0_0;
        end
        if(_zz_31) begin
          lruBit_10_0 <= _zz_lruBit_0_0;
        end
        if(_zz_32) begin
          lruBit_11_0 <= _zz_lruBit_0_0;
        end
        if(_zz_33) begin
          lruBit_12_0 <= _zz_lruBit_0_0;
        end
        if(_zz_34) begin
          lruBit_13_0 <= _zz_lruBit_0_0;
        end
        if(_zz_35) begin
          lruBit_14_0 <= _zz_lruBit_0_0;
        end
        if(_zz_36) begin
          lruBit_15_0 <= _zz_lruBit_0_0;
        end
        if(_zz_37) begin
          lruBit_16_0 <= _zz_lruBit_0_0;
        end
        if(_zz_38) begin
          lruBit_17_0 <= _zz_lruBit_0_0;
        end
        if(_zz_39) begin
          lruBit_18_0 <= _zz_lruBit_0_0;
        end
        if(_zz_40) begin
          lruBit_19_0 <= _zz_lruBit_0_0;
        end
        if(_zz_41) begin
          lruBit_20_0 <= _zz_lruBit_0_0;
        end
        if(_zz_42) begin
          lruBit_21_0 <= _zz_lruBit_0_0;
        end
        if(_zz_43) begin
          lruBit_22_0 <= _zz_lruBit_0_0;
        end
        if(_zz_44) begin
          lruBit_23_0 <= _zz_lruBit_0_0;
        end
        if(_zz_45) begin
          lruBit_24_0 <= _zz_lruBit_0_0;
        end
        if(_zz_46) begin
          lruBit_25_0 <= _zz_lruBit_0_0;
        end
        if(_zz_47) begin
          lruBit_26_0 <= _zz_lruBit_0_0;
        end
        if(_zz_48) begin
          lruBit_27_0 <= _zz_lruBit_0_0;
        end
        if(_zz_49) begin
          lruBit_28_0 <= _zz_lruBit_0_0;
        end
        if(_zz_50) begin
          lruBit_29_0 <= _zz_lruBit_0_0;
        end
        if(_zz_51) begin
          lruBit_30_0 <= _zz_lruBit_0_0;
        end
        if(_zz_52) begin
          lruBit_31_0 <= _zz_lruBit_0_0;
        end
        if(_zz_21) begin
          lruBit_0_1 <= _zz_lruBit_0_1;
        end
        if(_zz_22) begin
          lruBit_1_1 <= _zz_lruBit_0_1;
        end
        if(_zz_23) begin
          lruBit_2_1 <= _zz_lruBit_0_1;
        end
        if(_zz_24) begin
          lruBit_3_1 <= _zz_lruBit_0_1;
        end
        if(_zz_25) begin
          lruBit_4_1 <= _zz_lruBit_0_1;
        end
        if(_zz_26) begin
          lruBit_5_1 <= _zz_lruBit_0_1;
        end
        if(_zz_27) begin
          lruBit_6_1 <= _zz_lruBit_0_1;
        end
        if(_zz_28) begin
          lruBit_7_1 <= _zz_lruBit_0_1;
        end
        if(_zz_29) begin
          lruBit_8_1 <= _zz_lruBit_0_1;
        end
        if(_zz_30) begin
          lruBit_9_1 <= _zz_lruBit_0_1;
        end
        if(_zz_31) begin
          lruBit_10_1 <= _zz_lruBit_0_1;
        end
        if(_zz_32) begin
          lruBit_11_1 <= _zz_lruBit_0_1;
        end
        if(_zz_33) begin
          lruBit_12_1 <= _zz_lruBit_0_1;
        end
        if(_zz_34) begin
          lruBit_13_1 <= _zz_lruBit_0_1;
        end
        if(_zz_35) begin
          lruBit_14_1 <= _zz_lruBit_0_1;
        end
        if(_zz_36) begin
          lruBit_15_1 <= _zz_lruBit_0_1;
        end
        if(_zz_37) begin
          lruBit_16_1 <= _zz_lruBit_0_1;
        end
        if(_zz_38) begin
          lruBit_17_1 <= _zz_lruBit_0_1;
        end
        if(_zz_39) begin
          lruBit_18_1 <= _zz_lruBit_0_1;
        end
        if(_zz_40) begin
          lruBit_19_1 <= _zz_lruBit_0_1;
        end
        if(_zz_41) begin
          lruBit_20_1 <= _zz_lruBit_0_1;
        end
        if(_zz_42) begin
          lruBit_21_1 <= _zz_lruBit_0_1;
        end
        if(_zz_43) begin
          lruBit_22_1 <= _zz_lruBit_0_1;
        end
        if(_zz_44) begin
          lruBit_23_1 <= _zz_lruBit_0_1;
        end
        if(_zz_45) begin
          lruBit_24_1 <= _zz_lruBit_0_1;
        end
        if(_zz_46) begin
          lruBit_25_1 <= _zz_lruBit_0_1;
        end
        if(_zz_47) begin
          lruBit_26_1 <= _zz_lruBit_0_1;
        end
        if(_zz_48) begin
          lruBit_27_1 <= _zz_lruBit_0_1;
        end
        if(_zz_49) begin
          lruBit_28_1 <= _zz_lruBit_0_1;
        end
        if(_zz_50) begin
          lruBit_29_1 <= _zz_lruBit_0_1;
        end
        if(_zz_51) begin
          lruBit_30_1 <= _zz_lruBit_0_1;
        end
        if(_zz_52) begin
          lruBit_31_1 <= _zz_lruBit_0_1;
        end
        if(_zz_21) begin
          lruBit_0_2 <= _zz_lruBit_0_2;
        end
        if(_zz_22) begin
          lruBit_1_2 <= _zz_lruBit_0_2;
        end
        if(_zz_23) begin
          lruBit_2_2 <= _zz_lruBit_0_2;
        end
        if(_zz_24) begin
          lruBit_3_2 <= _zz_lruBit_0_2;
        end
        if(_zz_25) begin
          lruBit_4_2 <= _zz_lruBit_0_2;
        end
        if(_zz_26) begin
          lruBit_5_2 <= _zz_lruBit_0_2;
        end
        if(_zz_27) begin
          lruBit_6_2 <= _zz_lruBit_0_2;
        end
        if(_zz_28) begin
          lruBit_7_2 <= _zz_lruBit_0_2;
        end
        if(_zz_29) begin
          lruBit_8_2 <= _zz_lruBit_0_2;
        end
        if(_zz_30) begin
          lruBit_9_2 <= _zz_lruBit_0_2;
        end
        if(_zz_31) begin
          lruBit_10_2 <= _zz_lruBit_0_2;
        end
        if(_zz_32) begin
          lruBit_11_2 <= _zz_lruBit_0_2;
        end
        if(_zz_33) begin
          lruBit_12_2 <= _zz_lruBit_0_2;
        end
        if(_zz_34) begin
          lruBit_13_2 <= _zz_lruBit_0_2;
        end
        if(_zz_35) begin
          lruBit_14_2 <= _zz_lruBit_0_2;
        end
        if(_zz_36) begin
          lruBit_15_2 <= _zz_lruBit_0_2;
        end
        if(_zz_37) begin
          lruBit_16_2 <= _zz_lruBit_0_2;
        end
        if(_zz_38) begin
          lruBit_17_2 <= _zz_lruBit_0_2;
        end
        if(_zz_39) begin
          lruBit_18_2 <= _zz_lruBit_0_2;
        end
        if(_zz_40) begin
          lruBit_19_2 <= _zz_lruBit_0_2;
        end
        if(_zz_41) begin
          lruBit_20_2 <= _zz_lruBit_0_2;
        end
        if(_zz_42) begin
          lruBit_21_2 <= _zz_lruBit_0_2;
        end
        if(_zz_43) begin
          lruBit_22_2 <= _zz_lruBit_0_2;
        end
        if(_zz_44) begin
          lruBit_23_2 <= _zz_lruBit_0_2;
        end
        if(_zz_45) begin
          lruBit_24_2 <= _zz_lruBit_0_2;
        end
        if(_zz_46) begin
          lruBit_25_2 <= _zz_lruBit_0_2;
        end
        if(_zz_47) begin
          lruBit_26_2 <= _zz_lruBit_0_2;
        end
        if(_zz_48) begin
          lruBit_27_2 <= _zz_lruBit_0_2;
        end
        if(_zz_49) begin
          lruBit_28_2 <= _zz_lruBit_0_2;
        end
        if(_zz_50) begin
          lruBit_29_2 <= _zz_lruBit_0_2;
        end
        if(_zz_51) begin
          lruBit_30_2 <= _zz_lruBit_0_2;
        end
        if(_zz_52) begin
          lruBit_31_2 <= _zz_lruBit_0_2;
        end
      end
      if(dirtyUpdate) begin
        if(when_LSU_l341) begin
          if(_zz_53[0]) begin
            dirty_0_0 <= 1'b1;
          end
          if(_zz_53[1]) begin
            dirty_0_1 <= 1'b1;
          end
          if(_zz_53[2]) begin
            dirty_0_2 <= 1'b1;
          end
          if(_zz_53[3]) begin
            dirty_0_3 <= 1'b1;
          end
          if(_zz_53[4]) begin
            dirty_0_4 <= 1'b1;
          end
          if(_zz_53[5]) begin
            dirty_0_5 <= 1'b1;
          end
          if(_zz_53[6]) begin
            dirty_0_6 <= 1'b1;
          end
          if(_zz_53[7]) begin
            dirty_0_7 <= 1'b1;
          end
          if(_zz_53[8]) begin
            dirty_0_8 <= 1'b1;
          end
          if(_zz_53[9]) begin
            dirty_0_9 <= 1'b1;
          end
          if(_zz_53[10]) begin
            dirty_0_10 <= 1'b1;
          end
          if(_zz_53[11]) begin
            dirty_0_11 <= 1'b1;
          end
          if(_zz_53[12]) begin
            dirty_0_12 <= 1'b1;
          end
          if(_zz_53[13]) begin
            dirty_0_13 <= 1'b1;
          end
          if(_zz_53[14]) begin
            dirty_0_14 <= 1'b1;
          end
          if(_zz_53[15]) begin
            dirty_0_15 <= 1'b1;
          end
          if(_zz_53[16]) begin
            dirty_0_16 <= 1'b1;
          end
          if(_zz_53[17]) begin
            dirty_0_17 <= 1'b1;
          end
          if(_zz_53[18]) begin
            dirty_0_18 <= 1'b1;
          end
          if(_zz_53[19]) begin
            dirty_0_19 <= 1'b1;
          end
          if(_zz_53[20]) begin
            dirty_0_20 <= 1'b1;
          end
          if(_zz_53[21]) begin
            dirty_0_21 <= 1'b1;
          end
          if(_zz_53[22]) begin
            dirty_0_22 <= 1'b1;
          end
          if(_zz_53[23]) begin
            dirty_0_23 <= 1'b1;
          end
          if(_zz_53[24]) begin
            dirty_0_24 <= 1'b1;
          end
          if(_zz_53[25]) begin
            dirty_0_25 <= 1'b1;
          end
          if(_zz_53[26]) begin
            dirty_0_26 <= 1'b1;
          end
          if(_zz_53[27]) begin
            dirty_0_27 <= 1'b1;
          end
          if(_zz_53[28]) begin
            dirty_0_28 <= 1'b1;
          end
          if(_zz_53[29]) begin
            dirty_0_29 <= 1'b1;
          end
          if(_zz_53[30]) begin
            dirty_0_30 <= 1'b1;
          end
          if(_zz_53[31]) begin
            dirty_0_31 <= 1'b1;
          end
        end
        if(when_LSU_l341_1) begin
          if(_zz_54[0]) begin
            dirty_1_0 <= 1'b1;
          end
          if(_zz_54[1]) begin
            dirty_1_1 <= 1'b1;
          end
          if(_zz_54[2]) begin
            dirty_1_2 <= 1'b1;
          end
          if(_zz_54[3]) begin
            dirty_1_3 <= 1'b1;
          end
          if(_zz_54[4]) begin
            dirty_1_4 <= 1'b1;
          end
          if(_zz_54[5]) begin
            dirty_1_5 <= 1'b1;
          end
          if(_zz_54[6]) begin
            dirty_1_6 <= 1'b1;
          end
          if(_zz_54[7]) begin
            dirty_1_7 <= 1'b1;
          end
          if(_zz_54[8]) begin
            dirty_1_8 <= 1'b1;
          end
          if(_zz_54[9]) begin
            dirty_1_9 <= 1'b1;
          end
          if(_zz_54[10]) begin
            dirty_1_10 <= 1'b1;
          end
          if(_zz_54[11]) begin
            dirty_1_11 <= 1'b1;
          end
          if(_zz_54[12]) begin
            dirty_1_12 <= 1'b1;
          end
          if(_zz_54[13]) begin
            dirty_1_13 <= 1'b1;
          end
          if(_zz_54[14]) begin
            dirty_1_14 <= 1'b1;
          end
          if(_zz_54[15]) begin
            dirty_1_15 <= 1'b1;
          end
          if(_zz_54[16]) begin
            dirty_1_16 <= 1'b1;
          end
          if(_zz_54[17]) begin
            dirty_1_17 <= 1'b1;
          end
          if(_zz_54[18]) begin
            dirty_1_18 <= 1'b1;
          end
          if(_zz_54[19]) begin
            dirty_1_19 <= 1'b1;
          end
          if(_zz_54[20]) begin
            dirty_1_20 <= 1'b1;
          end
          if(_zz_54[21]) begin
            dirty_1_21 <= 1'b1;
          end
          if(_zz_54[22]) begin
            dirty_1_22 <= 1'b1;
          end
          if(_zz_54[23]) begin
            dirty_1_23 <= 1'b1;
          end
          if(_zz_54[24]) begin
            dirty_1_24 <= 1'b1;
          end
          if(_zz_54[25]) begin
            dirty_1_25 <= 1'b1;
          end
          if(_zz_54[26]) begin
            dirty_1_26 <= 1'b1;
          end
          if(_zz_54[27]) begin
            dirty_1_27 <= 1'b1;
          end
          if(_zz_54[28]) begin
            dirty_1_28 <= 1'b1;
          end
          if(_zz_54[29]) begin
            dirty_1_29 <= 1'b1;
          end
          if(_zz_54[30]) begin
            dirty_1_30 <= 1'b1;
          end
          if(_zz_54[31]) begin
            dirty_1_31 <= 1'b1;
          end
        end
        if(when_LSU_l341_2) begin
          if(_zz_55[0]) begin
            dirty_2_0 <= 1'b1;
          end
          if(_zz_55[1]) begin
            dirty_2_1 <= 1'b1;
          end
          if(_zz_55[2]) begin
            dirty_2_2 <= 1'b1;
          end
          if(_zz_55[3]) begin
            dirty_2_3 <= 1'b1;
          end
          if(_zz_55[4]) begin
            dirty_2_4 <= 1'b1;
          end
          if(_zz_55[5]) begin
            dirty_2_5 <= 1'b1;
          end
          if(_zz_55[6]) begin
            dirty_2_6 <= 1'b1;
          end
          if(_zz_55[7]) begin
            dirty_2_7 <= 1'b1;
          end
          if(_zz_55[8]) begin
            dirty_2_8 <= 1'b1;
          end
          if(_zz_55[9]) begin
            dirty_2_9 <= 1'b1;
          end
          if(_zz_55[10]) begin
            dirty_2_10 <= 1'b1;
          end
          if(_zz_55[11]) begin
            dirty_2_11 <= 1'b1;
          end
          if(_zz_55[12]) begin
            dirty_2_12 <= 1'b1;
          end
          if(_zz_55[13]) begin
            dirty_2_13 <= 1'b1;
          end
          if(_zz_55[14]) begin
            dirty_2_14 <= 1'b1;
          end
          if(_zz_55[15]) begin
            dirty_2_15 <= 1'b1;
          end
          if(_zz_55[16]) begin
            dirty_2_16 <= 1'b1;
          end
          if(_zz_55[17]) begin
            dirty_2_17 <= 1'b1;
          end
          if(_zz_55[18]) begin
            dirty_2_18 <= 1'b1;
          end
          if(_zz_55[19]) begin
            dirty_2_19 <= 1'b1;
          end
          if(_zz_55[20]) begin
            dirty_2_20 <= 1'b1;
          end
          if(_zz_55[21]) begin
            dirty_2_21 <= 1'b1;
          end
          if(_zz_55[22]) begin
            dirty_2_22 <= 1'b1;
          end
          if(_zz_55[23]) begin
            dirty_2_23 <= 1'b1;
          end
          if(_zz_55[24]) begin
            dirty_2_24 <= 1'b1;
          end
          if(_zz_55[25]) begin
            dirty_2_25 <= 1'b1;
          end
          if(_zz_55[26]) begin
            dirty_2_26 <= 1'b1;
          end
          if(_zz_55[27]) begin
            dirty_2_27 <= 1'b1;
          end
          if(_zz_55[28]) begin
            dirty_2_28 <= 1'b1;
          end
          if(_zz_55[29]) begin
            dirty_2_29 <= 1'b1;
          end
          if(_zz_55[30]) begin
            dirty_2_30 <= 1'b1;
          end
          if(_zz_55[31]) begin
            dirty_2_31 <= 1'b1;
          end
        end
        if(when_LSU_l341_3) begin
          if(_zz_56[0]) begin
            dirty_3_0 <= 1'b1;
          end
          if(_zz_56[1]) begin
            dirty_3_1 <= 1'b1;
          end
          if(_zz_56[2]) begin
            dirty_3_2 <= 1'b1;
          end
          if(_zz_56[3]) begin
            dirty_3_3 <= 1'b1;
          end
          if(_zz_56[4]) begin
            dirty_3_4 <= 1'b1;
          end
          if(_zz_56[5]) begin
            dirty_3_5 <= 1'b1;
          end
          if(_zz_56[6]) begin
            dirty_3_6 <= 1'b1;
          end
          if(_zz_56[7]) begin
            dirty_3_7 <= 1'b1;
          end
          if(_zz_56[8]) begin
            dirty_3_8 <= 1'b1;
          end
          if(_zz_56[9]) begin
            dirty_3_9 <= 1'b1;
          end
          if(_zz_56[10]) begin
            dirty_3_10 <= 1'b1;
          end
          if(_zz_56[11]) begin
            dirty_3_11 <= 1'b1;
          end
          if(_zz_56[12]) begin
            dirty_3_12 <= 1'b1;
          end
          if(_zz_56[13]) begin
            dirty_3_13 <= 1'b1;
          end
          if(_zz_56[14]) begin
            dirty_3_14 <= 1'b1;
          end
          if(_zz_56[15]) begin
            dirty_3_15 <= 1'b1;
          end
          if(_zz_56[16]) begin
            dirty_3_16 <= 1'b1;
          end
          if(_zz_56[17]) begin
            dirty_3_17 <= 1'b1;
          end
          if(_zz_56[18]) begin
            dirty_3_18 <= 1'b1;
          end
          if(_zz_56[19]) begin
            dirty_3_19 <= 1'b1;
          end
          if(_zz_56[20]) begin
            dirty_3_20 <= 1'b1;
          end
          if(_zz_56[21]) begin
            dirty_3_21 <= 1'b1;
          end
          if(_zz_56[22]) begin
            dirty_3_22 <= 1'b1;
          end
          if(_zz_56[23]) begin
            dirty_3_23 <= 1'b1;
          end
          if(_zz_56[24]) begin
            dirty_3_24 <= 1'b1;
          end
          if(_zz_56[25]) begin
            dirty_3_25 <= 1'b1;
          end
          if(_zz_56[26]) begin
            dirty_3_26 <= 1'b1;
          end
          if(_zz_56[27]) begin
            dirty_3_27 <= 1'b1;
          end
          if(_zz_56[28]) begin
            dirty_3_28 <= 1'b1;
          end
          if(_zz_56[29]) begin
            dirty_3_29 <= 1'b1;
          end
          if(_zz_56[30]) begin
            dirty_3_30 <= 1'b1;
          end
          if(_zz_56[31]) begin
            dirty_3_31 <= 1'b1;
          end
        end
      end
      if(refilling) begin
        if(when_LSU_l348) begin
          if(_zz_57[0]) begin
            dirty_0_0 <= latestWrite_prevDirty;
          end
          if(_zz_57[1]) begin
            dirty_0_1 <= latestWrite_prevDirty;
          end
          if(_zz_57[2]) begin
            dirty_0_2 <= latestWrite_prevDirty;
          end
          if(_zz_57[3]) begin
            dirty_0_3 <= latestWrite_prevDirty;
          end
          if(_zz_57[4]) begin
            dirty_0_4 <= latestWrite_prevDirty;
          end
          if(_zz_57[5]) begin
            dirty_0_5 <= latestWrite_prevDirty;
          end
          if(_zz_57[6]) begin
            dirty_0_6 <= latestWrite_prevDirty;
          end
          if(_zz_57[7]) begin
            dirty_0_7 <= latestWrite_prevDirty;
          end
          if(_zz_57[8]) begin
            dirty_0_8 <= latestWrite_prevDirty;
          end
          if(_zz_57[9]) begin
            dirty_0_9 <= latestWrite_prevDirty;
          end
          if(_zz_57[10]) begin
            dirty_0_10 <= latestWrite_prevDirty;
          end
          if(_zz_57[11]) begin
            dirty_0_11 <= latestWrite_prevDirty;
          end
          if(_zz_57[12]) begin
            dirty_0_12 <= latestWrite_prevDirty;
          end
          if(_zz_57[13]) begin
            dirty_0_13 <= latestWrite_prevDirty;
          end
          if(_zz_57[14]) begin
            dirty_0_14 <= latestWrite_prevDirty;
          end
          if(_zz_57[15]) begin
            dirty_0_15 <= latestWrite_prevDirty;
          end
          if(_zz_57[16]) begin
            dirty_0_16 <= latestWrite_prevDirty;
          end
          if(_zz_57[17]) begin
            dirty_0_17 <= latestWrite_prevDirty;
          end
          if(_zz_57[18]) begin
            dirty_0_18 <= latestWrite_prevDirty;
          end
          if(_zz_57[19]) begin
            dirty_0_19 <= latestWrite_prevDirty;
          end
          if(_zz_57[20]) begin
            dirty_0_20 <= latestWrite_prevDirty;
          end
          if(_zz_57[21]) begin
            dirty_0_21 <= latestWrite_prevDirty;
          end
          if(_zz_57[22]) begin
            dirty_0_22 <= latestWrite_prevDirty;
          end
          if(_zz_57[23]) begin
            dirty_0_23 <= latestWrite_prevDirty;
          end
          if(_zz_57[24]) begin
            dirty_0_24 <= latestWrite_prevDirty;
          end
          if(_zz_57[25]) begin
            dirty_0_25 <= latestWrite_prevDirty;
          end
          if(_zz_57[26]) begin
            dirty_0_26 <= latestWrite_prevDirty;
          end
          if(_zz_57[27]) begin
            dirty_0_27 <= latestWrite_prevDirty;
          end
          if(_zz_57[28]) begin
            dirty_0_28 <= latestWrite_prevDirty;
          end
          if(_zz_57[29]) begin
            dirty_0_29 <= latestWrite_prevDirty;
          end
          if(_zz_57[30]) begin
            dirty_0_30 <= latestWrite_prevDirty;
          end
          if(_zz_57[31]) begin
            dirty_0_31 <= latestWrite_prevDirty;
          end
        end
        if(when_LSU_l348_1) begin
          if(_zz_58[0]) begin
            dirty_1_0 <= latestWrite_prevDirty;
          end
          if(_zz_58[1]) begin
            dirty_1_1 <= latestWrite_prevDirty;
          end
          if(_zz_58[2]) begin
            dirty_1_2 <= latestWrite_prevDirty;
          end
          if(_zz_58[3]) begin
            dirty_1_3 <= latestWrite_prevDirty;
          end
          if(_zz_58[4]) begin
            dirty_1_4 <= latestWrite_prevDirty;
          end
          if(_zz_58[5]) begin
            dirty_1_5 <= latestWrite_prevDirty;
          end
          if(_zz_58[6]) begin
            dirty_1_6 <= latestWrite_prevDirty;
          end
          if(_zz_58[7]) begin
            dirty_1_7 <= latestWrite_prevDirty;
          end
          if(_zz_58[8]) begin
            dirty_1_8 <= latestWrite_prevDirty;
          end
          if(_zz_58[9]) begin
            dirty_1_9 <= latestWrite_prevDirty;
          end
          if(_zz_58[10]) begin
            dirty_1_10 <= latestWrite_prevDirty;
          end
          if(_zz_58[11]) begin
            dirty_1_11 <= latestWrite_prevDirty;
          end
          if(_zz_58[12]) begin
            dirty_1_12 <= latestWrite_prevDirty;
          end
          if(_zz_58[13]) begin
            dirty_1_13 <= latestWrite_prevDirty;
          end
          if(_zz_58[14]) begin
            dirty_1_14 <= latestWrite_prevDirty;
          end
          if(_zz_58[15]) begin
            dirty_1_15 <= latestWrite_prevDirty;
          end
          if(_zz_58[16]) begin
            dirty_1_16 <= latestWrite_prevDirty;
          end
          if(_zz_58[17]) begin
            dirty_1_17 <= latestWrite_prevDirty;
          end
          if(_zz_58[18]) begin
            dirty_1_18 <= latestWrite_prevDirty;
          end
          if(_zz_58[19]) begin
            dirty_1_19 <= latestWrite_prevDirty;
          end
          if(_zz_58[20]) begin
            dirty_1_20 <= latestWrite_prevDirty;
          end
          if(_zz_58[21]) begin
            dirty_1_21 <= latestWrite_prevDirty;
          end
          if(_zz_58[22]) begin
            dirty_1_22 <= latestWrite_prevDirty;
          end
          if(_zz_58[23]) begin
            dirty_1_23 <= latestWrite_prevDirty;
          end
          if(_zz_58[24]) begin
            dirty_1_24 <= latestWrite_prevDirty;
          end
          if(_zz_58[25]) begin
            dirty_1_25 <= latestWrite_prevDirty;
          end
          if(_zz_58[26]) begin
            dirty_1_26 <= latestWrite_prevDirty;
          end
          if(_zz_58[27]) begin
            dirty_1_27 <= latestWrite_prevDirty;
          end
          if(_zz_58[28]) begin
            dirty_1_28 <= latestWrite_prevDirty;
          end
          if(_zz_58[29]) begin
            dirty_1_29 <= latestWrite_prevDirty;
          end
          if(_zz_58[30]) begin
            dirty_1_30 <= latestWrite_prevDirty;
          end
          if(_zz_58[31]) begin
            dirty_1_31 <= latestWrite_prevDirty;
          end
        end
        if(when_LSU_l348_2) begin
          if(_zz_59[0]) begin
            dirty_2_0 <= latestWrite_prevDirty;
          end
          if(_zz_59[1]) begin
            dirty_2_1 <= latestWrite_prevDirty;
          end
          if(_zz_59[2]) begin
            dirty_2_2 <= latestWrite_prevDirty;
          end
          if(_zz_59[3]) begin
            dirty_2_3 <= latestWrite_prevDirty;
          end
          if(_zz_59[4]) begin
            dirty_2_4 <= latestWrite_prevDirty;
          end
          if(_zz_59[5]) begin
            dirty_2_5 <= latestWrite_prevDirty;
          end
          if(_zz_59[6]) begin
            dirty_2_6 <= latestWrite_prevDirty;
          end
          if(_zz_59[7]) begin
            dirty_2_7 <= latestWrite_prevDirty;
          end
          if(_zz_59[8]) begin
            dirty_2_8 <= latestWrite_prevDirty;
          end
          if(_zz_59[9]) begin
            dirty_2_9 <= latestWrite_prevDirty;
          end
          if(_zz_59[10]) begin
            dirty_2_10 <= latestWrite_prevDirty;
          end
          if(_zz_59[11]) begin
            dirty_2_11 <= latestWrite_prevDirty;
          end
          if(_zz_59[12]) begin
            dirty_2_12 <= latestWrite_prevDirty;
          end
          if(_zz_59[13]) begin
            dirty_2_13 <= latestWrite_prevDirty;
          end
          if(_zz_59[14]) begin
            dirty_2_14 <= latestWrite_prevDirty;
          end
          if(_zz_59[15]) begin
            dirty_2_15 <= latestWrite_prevDirty;
          end
          if(_zz_59[16]) begin
            dirty_2_16 <= latestWrite_prevDirty;
          end
          if(_zz_59[17]) begin
            dirty_2_17 <= latestWrite_prevDirty;
          end
          if(_zz_59[18]) begin
            dirty_2_18 <= latestWrite_prevDirty;
          end
          if(_zz_59[19]) begin
            dirty_2_19 <= latestWrite_prevDirty;
          end
          if(_zz_59[20]) begin
            dirty_2_20 <= latestWrite_prevDirty;
          end
          if(_zz_59[21]) begin
            dirty_2_21 <= latestWrite_prevDirty;
          end
          if(_zz_59[22]) begin
            dirty_2_22 <= latestWrite_prevDirty;
          end
          if(_zz_59[23]) begin
            dirty_2_23 <= latestWrite_prevDirty;
          end
          if(_zz_59[24]) begin
            dirty_2_24 <= latestWrite_prevDirty;
          end
          if(_zz_59[25]) begin
            dirty_2_25 <= latestWrite_prevDirty;
          end
          if(_zz_59[26]) begin
            dirty_2_26 <= latestWrite_prevDirty;
          end
          if(_zz_59[27]) begin
            dirty_2_27 <= latestWrite_prevDirty;
          end
          if(_zz_59[28]) begin
            dirty_2_28 <= latestWrite_prevDirty;
          end
          if(_zz_59[29]) begin
            dirty_2_29 <= latestWrite_prevDirty;
          end
          if(_zz_59[30]) begin
            dirty_2_30 <= latestWrite_prevDirty;
          end
          if(_zz_59[31]) begin
            dirty_2_31 <= latestWrite_prevDirty;
          end
        end
        if(when_LSU_l348_3) begin
          if(_zz_60[0]) begin
            dirty_3_0 <= latestWrite_prevDirty;
          end
          if(_zz_60[1]) begin
            dirty_3_1 <= latestWrite_prevDirty;
          end
          if(_zz_60[2]) begin
            dirty_3_2 <= latestWrite_prevDirty;
          end
          if(_zz_60[3]) begin
            dirty_3_3 <= latestWrite_prevDirty;
          end
          if(_zz_60[4]) begin
            dirty_3_4 <= latestWrite_prevDirty;
          end
          if(_zz_60[5]) begin
            dirty_3_5 <= latestWrite_prevDirty;
          end
          if(_zz_60[6]) begin
            dirty_3_6 <= latestWrite_prevDirty;
          end
          if(_zz_60[7]) begin
            dirty_3_7 <= latestWrite_prevDirty;
          end
          if(_zz_60[8]) begin
            dirty_3_8 <= latestWrite_prevDirty;
          end
          if(_zz_60[9]) begin
            dirty_3_9 <= latestWrite_prevDirty;
          end
          if(_zz_60[10]) begin
            dirty_3_10 <= latestWrite_prevDirty;
          end
          if(_zz_60[11]) begin
            dirty_3_11 <= latestWrite_prevDirty;
          end
          if(_zz_60[12]) begin
            dirty_3_12 <= latestWrite_prevDirty;
          end
          if(_zz_60[13]) begin
            dirty_3_13 <= latestWrite_prevDirty;
          end
          if(_zz_60[14]) begin
            dirty_3_14 <= latestWrite_prevDirty;
          end
          if(_zz_60[15]) begin
            dirty_3_15 <= latestWrite_prevDirty;
          end
          if(_zz_60[16]) begin
            dirty_3_16 <= latestWrite_prevDirty;
          end
          if(_zz_60[17]) begin
            dirty_3_17 <= latestWrite_prevDirty;
          end
          if(_zz_60[18]) begin
            dirty_3_18 <= latestWrite_prevDirty;
          end
          if(_zz_60[19]) begin
            dirty_3_19 <= latestWrite_prevDirty;
          end
          if(_zz_60[20]) begin
            dirty_3_20 <= latestWrite_prevDirty;
          end
          if(_zz_60[21]) begin
            dirty_3_21 <= latestWrite_prevDirty;
          end
          if(_zz_60[22]) begin
            dirty_3_22 <= latestWrite_prevDirty;
          end
          if(_zz_60[23]) begin
            dirty_3_23 <= latestWrite_prevDirty;
          end
          if(_zz_60[24]) begin
            dirty_3_24 <= latestWrite_prevDirty;
          end
          if(_zz_60[25]) begin
            dirty_3_25 <= latestWrite_prevDirty;
          end
          if(_zz_60[26]) begin
            dirty_3_26 <= latestWrite_prevDirty;
          end
          if(_zz_60[27]) begin
            dirty_3_27 <= latestWrite_prevDirty;
          end
          if(_zz_60[28]) begin
            dirty_3_28 <= latestWrite_prevDirty;
          end
          if(_zz_60[29]) begin
            dirty_3_29 <= latestWrite_prevDirty;
          end
          if(_zz_60[30]) begin
            dirty_3_30 <= latestWrite_prevDirty;
          end
          if(_zz_60[31]) begin
            dirty_3_31 <= latestWrite_prevDirty;
          end
        end
      end
      if(stage1Out_fire) begin
        if(when_LSU_l357) begin
          wayDirtyBypass <= (axiLoad ? transferWaySelect : hit);
        end else begin
          wayDirtyBypass <= 4'b0000;
        end
      end
      if(when_LSU_l661) begin
        if(when_LSU_l663) begin
          if(_zz_61[0]) begin
            valid_0_0 <= 1'b0;
          end
          if(_zz_61[1]) begin
            valid_0_1 <= 1'b0;
          end
          if(_zz_61[2]) begin
            valid_0_2 <= 1'b0;
          end
          if(_zz_61[3]) begin
            valid_0_3 <= 1'b0;
          end
          if(_zz_61[4]) begin
            valid_0_4 <= 1'b0;
          end
          if(_zz_61[5]) begin
            valid_0_5 <= 1'b0;
          end
          if(_zz_61[6]) begin
            valid_0_6 <= 1'b0;
          end
          if(_zz_61[7]) begin
            valid_0_7 <= 1'b0;
          end
          if(_zz_61[8]) begin
            valid_0_8 <= 1'b0;
          end
          if(_zz_61[9]) begin
            valid_0_9 <= 1'b0;
          end
          if(_zz_61[10]) begin
            valid_0_10 <= 1'b0;
          end
          if(_zz_61[11]) begin
            valid_0_11 <= 1'b0;
          end
          if(_zz_61[12]) begin
            valid_0_12 <= 1'b0;
          end
          if(_zz_61[13]) begin
            valid_0_13 <= 1'b0;
          end
          if(_zz_61[14]) begin
            valid_0_14 <= 1'b0;
          end
          if(_zz_61[15]) begin
            valid_0_15 <= 1'b0;
          end
          if(_zz_61[16]) begin
            valid_0_16 <= 1'b0;
          end
          if(_zz_61[17]) begin
            valid_0_17 <= 1'b0;
          end
          if(_zz_61[18]) begin
            valid_0_18 <= 1'b0;
          end
          if(_zz_61[19]) begin
            valid_0_19 <= 1'b0;
          end
          if(_zz_61[20]) begin
            valid_0_20 <= 1'b0;
          end
          if(_zz_61[21]) begin
            valid_0_21 <= 1'b0;
          end
          if(_zz_61[22]) begin
            valid_0_22 <= 1'b0;
          end
          if(_zz_61[23]) begin
            valid_0_23 <= 1'b0;
          end
          if(_zz_61[24]) begin
            valid_0_24 <= 1'b0;
          end
          if(_zz_61[25]) begin
            valid_0_25 <= 1'b0;
          end
          if(_zz_61[26]) begin
            valid_0_26 <= 1'b0;
          end
          if(_zz_61[27]) begin
            valid_0_27 <= 1'b0;
          end
          if(_zz_61[28]) begin
            valid_0_28 <= 1'b0;
          end
          if(_zz_61[29]) begin
            valid_0_29 <= 1'b0;
          end
          if(_zz_61[30]) begin
            valid_0_30 <= 1'b0;
          end
          if(_zz_61[31]) begin
            valid_0_31 <= 1'b0;
          end
        end
        if(when_LSU_l663_1) begin
          if(_zz_62[0]) begin
            valid_1_0 <= 1'b0;
          end
          if(_zz_62[1]) begin
            valid_1_1 <= 1'b0;
          end
          if(_zz_62[2]) begin
            valid_1_2 <= 1'b0;
          end
          if(_zz_62[3]) begin
            valid_1_3 <= 1'b0;
          end
          if(_zz_62[4]) begin
            valid_1_4 <= 1'b0;
          end
          if(_zz_62[5]) begin
            valid_1_5 <= 1'b0;
          end
          if(_zz_62[6]) begin
            valid_1_6 <= 1'b0;
          end
          if(_zz_62[7]) begin
            valid_1_7 <= 1'b0;
          end
          if(_zz_62[8]) begin
            valid_1_8 <= 1'b0;
          end
          if(_zz_62[9]) begin
            valid_1_9 <= 1'b0;
          end
          if(_zz_62[10]) begin
            valid_1_10 <= 1'b0;
          end
          if(_zz_62[11]) begin
            valid_1_11 <= 1'b0;
          end
          if(_zz_62[12]) begin
            valid_1_12 <= 1'b0;
          end
          if(_zz_62[13]) begin
            valid_1_13 <= 1'b0;
          end
          if(_zz_62[14]) begin
            valid_1_14 <= 1'b0;
          end
          if(_zz_62[15]) begin
            valid_1_15 <= 1'b0;
          end
          if(_zz_62[16]) begin
            valid_1_16 <= 1'b0;
          end
          if(_zz_62[17]) begin
            valid_1_17 <= 1'b0;
          end
          if(_zz_62[18]) begin
            valid_1_18 <= 1'b0;
          end
          if(_zz_62[19]) begin
            valid_1_19 <= 1'b0;
          end
          if(_zz_62[20]) begin
            valid_1_20 <= 1'b0;
          end
          if(_zz_62[21]) begin
            valid_1_21 <= 1'b0;
          end
          if(_zz_62[22]) begin
            valid_1_22 <= 1'b0;
          end
          if(_zz_62[23]) begin
            valid_1_23 <= 1'b0;
          end
          if(_zz_62[24]) begin
            valid_1_24 <= 1'b0;
          end
          if(_zz_62[25]) begin
            valid_1_25 <= 1'b0;
          end
          if(_zz_62[26]) begin
            valid_1_26 <= 1'b0;
          end
          if(_zz_62[27]) begin
            valid_1_27 <= 1'b0;
          end
          if(_zz_62[28]) begin
            valid_1_28 <= 1'b0;
          end
          if(_zz_62[29]) begin
            valid_1_29 <= 1'b0;
          end
          if(_zz_62[30]) begin
            valid_1_30 <= 1'b0;
          end
          if(_zz_62[31]) begin
            valid_1_31 <= 1'b0;
          end
        end
        if(when_LSU_l663_2) begin
          if(_zz_63[0]) begin
            valid_2_0 <= 1'b0;
          end
          if(_zz_63[1]) begin
            valid_2_1 <= 1'b0;
          end
          if(_zz_63[2]) begin
            valid_2_2 <= 1'b0;
          end
          if(_zz_63[3]) begin
            valid_2_3 <= 1'b0;
          end
          if(_zz_63[4]) begin
            valid_2_4 <= 1'b0;
          end
          if(_zz_63[5]) begin
            valid_2_5 <= 1'b0;
          end
          if(_zz_63[6]) begin
            valid_2_6 <= 1'b0;
          end
          if(_zz_63[7]) begin
            valid_2_7 <= 1'b0;
          end
          if(_zz_63[8]) begin
            valid_2_8 <= 1'b0;
          end
          if(_zz_63[9]) begin
            valid_2_9 <= 1'b0;
          end
          if(_zz_63[10]) begin
            valid_2_10 <= 1'b0;
          end
          if(_zz_63[11]) begin
            valid_2_11 <= 1'b0;
          end
          if(_zz_63[12]) begin
            valid_2_12 <= 1'b0;
          end
          if(_zz_63[13]) begin
            valid_2_13 <= 1'b0;
          end
          if(_zz_63[14]) begin
            valid_2_14 <= 1'b0;
          end
          if(_zz_63[15]) begin
            valid_2_15 <= 1'b0;
          end
          if(_zz_63[16]) begin
            valid_2_16 <= 1'b0;
          end
          if(_zz_63[17]) begin
            valid_2_17 <= 1'b0;
          end
          if(_zz_63[18]) begin
            valid_2_18 <= 1'b0;
          end
          if(_zz_63[19]) begin
            valid_2_19 <= 1'b0;
          end
          if(_zz_63[20]) begin
            valid_2_20 <= 1'b0;
          end
          if(_zz_63[21]) begin
            valid_2_21 <= 1'b0;
          end
          if(_zz_63[22]) begin
            valid_2_22 <= 1'b0;
          end
          if(_zz_63[23]) begin
            valid_2_23 <= 1'b0;
          end
          if(_zz_63[24]) begin
            valid_2_24 <= 1'b0;
          end
          if(_zz_63[25]) begin
            valid_2_25 <= 1'b0;
          end
          if(_zz_63[26]) begin
            valid_2_26 <= 1'b0;
          end
          if(_zz_63[27]) begin
            valid_2_27 <= 1'b0;
          end
          if(_zz_63[28]) begin
            valid_2_28 <= 1'b0;
          end
          if(_zz_63[29]) begin
            valid_2_29 <= 1'b0;
          end
          if(_zz_63[30]) begin
            valid_2_30 <= 1'b0;
          end
          if(_zz_63[31]) begin
            valid_2_31 <= 1'b0;
          end
        end
        if(when_LSU_l663_3) begin
          if(_zz_64[0]) begin
            valid_3_0 <= 1'b0;
          end
          if(_zz_64[1]) begin
            valid_3_1 <= 1'b0;
          end
          if(_zz_64[2]) begin
            valid_3_2 <= 1'b0;
          end
          if(_zz_64[3]) begin
            valid_3_3 <= 1'b0;
          end
          if(_zz_64[4]) begin
            valid_3_4 <= 1'b0;
          end
          if(_zz_64[5]) begin
            valid_3_5 <= 1'b0;
          end
          if(_zz_64[6]) begin
            valid_3_6 <= 1'b0;
          end
          if(_zz_64[7]) begin
            valid_3_7 <= 1'b0;
          end
          if(_zz_64[8]) begin
            valid_3_8 <= 1'b0;
          end
          if(_zz_64[9]) begin
            valid_3_9 <= 1'b0;
          end
          if(_zz_64[10]) begin
            valid_3_10 <= 1'b0;
          end
          if(_zz_64[11]) begin
            valid_3_11 <= 1'b0;
          end
          if(_zz_64[12]) begin
            valid_3_12 <= 1'b0;
          end
          if(_zz_64[13]) begin
            valid_3_13 <= 1'b0;
          end
          if(_zz_64[14]) begin
            valid_3_14 <= 1'b0;
          end
          if(_zz_64[15]) begin
            valid_3_15 <= 1'b0;
          end
          if(_zz_64[16]) begin
            valid_3_16 <= 1'b0;
          end
          if(_zz_64[17]) begin
            valid_3_17 <= 1'b0;
          end
          if(_zz_64[18]) begin
            valid_3_18 <= 1'b0;
          end
          if(_zz_64[19]) begin
            valid_3_19 <= 1'b0;
          end
          if(_zz_64[20]) begin
            valid_3_20 <= 1'b0;
          end
          if(_zz_64[21]) begin
            valid_3_21 <= 1'b0;
          end
          if(_zz_64[22]) begin
            valid_3_22 <= 1'b0;
          end
          if(_zz_64[23]) begin
            valid_3_23 <= 1'b0;
          end
          if(_zz_64[24]) begin
            valid_3_24 <= 1'b0;
          end
          if(_zz_64[25]) begin
            valid_3_25 <= 1'b0;
          end
          if(_zz_64[26]) begin
            valid_3_26 <= 1'b0;
          end
          if(_zz_64[27]) begin
            valid_3_27 <= 1'b0;
          end
          if(_zz_64[28]) begin
            valid_3_28 <= 1'b0;
          end
          if(_zz_64[29]) begin
            valid_3_29 <= 1'b0;
          end
          if(_zz_64[30]) begin
            valid_3_30 <= 1'b0;
          end
          if(_zz_64[31]) begin
            valid_3_31 <= 1'b0;
          end
        end
      end
      axiCtrl_stateReg <= axiCtrl_stateNext;
      case(axiCtrl_stateReg)
        axiCtrl_enumDef_idle : begin
          if(when_LSU_l436) begin
            transferRAddrHi <= missingEntry_paddr[31 : 6];
            transferRAddrMid <= missingEntry_paddr[5 : 2];
            transferRAddrLo <= missingEntry_paddr[1 : 0];
            transferWAddrHi <= (missingEntry_uncached ? missingEntry_paddr[31 : 6] : missingEntry_prevPaddr[31 : 6]);
            transferWAddrMid <= (missingEntry_uncached ? missingEntry_paddr[5 : 2] : 4'b0000);
            transferWAddrLo <= (missingEntry_uncached ? missingEntry_paddr[1 : 0] : 2'b00);
            transferUncached <= missingEntry_uncached;
            transferWaySelect <= missingEntry_waySelect;
            transferWData <= missingEntry_storeData;
            transferLSMask <= missingEntry_lsMask;
          end
          if(when_LSU_l453) begin
            transferWAddrHi <= cacopPAddr[31 : 6];
            transferWAddrMid <= cacopPAddr[5 : 2];
            transferWAddrLo <= cacopPAddr[1 : 0];
            transferCACOP <= 1'b1;
            transferUncached <= 1'b0;
            transferWaySelect <= cacopWay;
          end
        end
        axiCtrl_enumDef_readReq : begin
          if(when_LSU_l471) begin
            if(when_LSU_l473) begin
              if(_zz_65[0]) begin
                valid_0_0 <= 1'b1;
              end
              if(_zz_65[1]) begin
                valid_0_1 <= 1'b1;
              end
              if(_zz_65[2]) begin
                valid_0_2 <= 1'b1;
              end
              if(_zz_65[3]) begin
                valid_0_3 <= 1'b1;
              end
              if(_zz_65[4]) begin
                valid_0_4 <= 1'b1;
              end
              if(_zz_65[5]) begin
                valid_0_5 <= 1'b1;
              end
              if(_zz_65[6]) begin
                valid_0_6 <= 1'b1;
              end
              if(_zz_65[7]) begin
                valid_0_7 <= 1'b1;
              end
              if(_zz_65[8]) begin
                valid_0_8 <= 1'b1;
              end
              if(_zz_65[9]) begin
                valid_0_9 <= 1'b1;
              end
              if(_zz_65[10]) begin
                valid_0_10 <= 1'b1;
              end
              if(_zz_65[11]) begin
                valid_0_11 <= 1'b1;
              end
              if(_zz_65[12]) begin
                valid_0_12 <= 1'b1;
              end
              if(_zz_65[13]) begin
                valid_0_13 <= 1'b1;
              end
              if(_zz_65[14]) begin
                valid_0_14 <= 1'b1;
              end
              if(_zz_65[15]) begin
                valid_0_15 <= 1'b1;
              end
              if(_zz_65[16]) begin
                valid_0_16 <= 1'b1;
              end
              if(_zz_65[17]) begin
                valid_0_17 <= 1'b1;
              end
              if(_zz_65[18]) begin
                valid_0_18 <= 1'b1;
              end
              if(_zz_65[19]) begin
                valid_0_19 <= 1'b1;
              end
              if(_zz_65[20]) begin
                valid_0_20 <= 1'b1;
              end
              if(_zz_65[21]) begin
                valid_0_21 <= 1'b1;
              end
              if(_zz_65[22]) begin
                valid_0_22 <= 1'b1;
              end
              if(_zz_65[23]) begin
                valid_0_23 <= 1'b1;
              end
              if(_zz_65[24]) begin
                valid_0_24 <= 1'b1;
              end
              if(_zz_65[25]) begin
                valid_0_25 <= 1'b1;
              end
              if(_zz_65[26]) begin
                valid_0_26 <= 1'b1;
              end
              if(_zz_65[27]) begin
                valid_0_27 <= 1'b1;
              end
              if(_zz_65[28]) begin
                valid_0_28 <= 1'b1;
              end
              if(_zz_65[29]) begin
                valid_0_29 <= 1'b1;
              end
              if(_zz_65[30]) begin
                valid_0_30 <= 1'b1;
              end
              if(_zz_65[31]) begin
                valid_0_31 <= 1'b1;
              end
              if(_zz_66[0]) begin
                dirty_0_0 <= 1'b0;
              end
              if(_zz_66[1]) begin
                dirty_0_1 <= 1'b0;
              end
              if(_zz_66[2]) begin
                dirty_0_2 <= 1'b0;
              end
              if(_zz_66[3]) begin
                dirty_0_3 <= 1'b0;
              end
              if(_zz_66[4]) begin
                dirty_0_4 <= 1'b0;
              end
              if(_zz_66[5]) begin
                dirty_0_5 <= 1'b0;
              end
              if(_zz_66[6]) begin
                dirty_0_6 <= 1'b0;
              end
              if(_zz_66[7]) begin
                dirty_0_7 <= 1'b0;
              end
              if(_zz_66[8]) begin
                dirty_0_8 <= 1'b0;
              end
              if(_zz_66[9]) begin
                dirty_0_9 <= 1'b0;
              end
              if(_zz_66[10]) begin
                dirty_0_10 <= 1'b0;
              end
              if(_zz_66[11]) begin
                dirty_0_11 <= 1'b0;
              end
              if(_zz_66[12]) begin
                dirty_0_12 <= 1'b0;
              end
              if(_zz_66[13]) begin
                dirty_0_13 <= 1'b0;
              end
              if(_zz_66[14]) begin
                dirty_0_14 <= 1'b0;
              end
              if(_zz_66[15]) begin
                dirty_0_15 <= 1'b0;
              end
              if(_zz_66[16]) begin
                dirty_0_16 <= 1'b0;
              end
              if(_zz_66[17]) begin
                dirty_0_17 <= 1'b0;
              end
              if(_zz_66[18]) begin
                dirty_0_18 <= 1'b0;
              end
              if(_zz_66[19]) begin
                dirty_0_19 <= 1'b0;
              end
              if(_zz_66[20]) begin
                dirty_0_20 <= 1'b0;
              end
              if(_zz_66[21]) begin
                dirty_0_21 <= 1'b0;
              end
              if(_zz_66[22]) begin
                dirty_0_22 <= 1'b0;
              end
              if(_zz_66[23]) begin
                dirty_0_23 <= 1'b0;
              end
              if(_zz_66[24]) begin
                dirty_0_24 <= 1'b0;
              end
              if(_zz_66[25]) begin
                dirty_0_25 <= 1'b0;
              end
              if(_zz_66[26]) begin
                dirty_0_26 <= 1'b0;
              end
              if(_zz_66[27]) begin
                dirty_0_27 <= 1'b0;
              end
              if(_zz_66[28]) begin
                dirty_0_28 <= 1'b0;
              end
              if(_zz_66[29]) begin
                dirty_0_29 <= 1'b0;
              end
              if(_zz_66[30]) begin
                dirty_0_30 <= 1'b0;
              end
              if(_zz_66[31]) begin
                dirty_0_31 <= 1'b0;
              end
            end
            if(when_LSU_l473_1) begin
              if(_zz_67[0]) begin
                valid_1_0 <= 1'b1;
              end
              if(_zz_67[1]) begin
                valid_1_1 <= 1'b1;
              end
              if(_zz_67[2]) begin
                valid_1_2 <= 1'b1;
              end
              if(_zz_67[3]) begin
                valid_1_3 <= 1'b1;
              end
              if(_zz_67[4]) begin
                valid_1_4 <= 1'b1;
              end
              if(_zz_67[5]) begin
                valid_1_5 <= 1'b1;
              end
              if(_zz_67[6]) begin
                valid_1_6 <= 1'b1;
              end
              if(_zz_67[7]) begin
                valid_1_7 <= 1'b1;
              end
              if(_zz_67[8]) begin
                valid_1_8 <= 1'b1;
              end
              if(_zz_67[9]) begin
                valid_1_9 <= 1'b1;
              end
              if(_zz_67[10]) begin
                valid_1_10 <= 1'b1;
              end
              if(_zz_67[11]) begin
                valid_1_11 <= 1'b1;
              end
              if(_zz_67[12]) begin
                valid_1_12 <= 1'b1;
              end
              if(_zz_67[13]) begin
                valid_1_13 <= 1'b1;
              end
              if(_zz_67[14]) begin
                valid_1_14 <= 1'b1;
              end
              if(_zz_67[15]) begin
                valid_1_15 <= 1'b1;
              end
              if(_zz_67[16]) begin
                valid_1_16 <= 1'b1;
              end
              if(_zz_67[17]) begin
                valid_1_17 <= 1'b1;
              end
              if(_zz_67[18]) begin
                valid_1_18 <= 1'b1;
              end
              if(_zz_67[19]) begin
                valid_1_19 <= 1'b1;
              end
              if(_zz_67[20]) begin
                valid_1_20 <= 1'b1;
              end
              if(_zz_67[21]) begin
                valid_1_21 <= 1'b1;
              end
              if(_zz_67[22]) begin
                valid_1_22 <= 1'b1;
              end
              if(_zz_67[23]) begin
                valid_1_23 <= 1'b1;
              end
              if(_zz_67[24]) begin
                valid_1_24 <= 1'b1;
              end
              if(_zz_67[25]) begin
                valid_1_25 <= 1'b1;
              end
              if(_zz_67[26]) begin
                valid_1_26 <= 1'b1;
              end
              if(_zz_67[27]) begin
                valid_1_27 <= 1'b1;
              end
              if(_zz_67[28]) begin
                valid_1_28 <= 1'b1;
              end
              if(_zz_67[29]) begin
                valid_1_29 <= 1'b1;
              end
              if(_zz_67[30]) begin
                valid_1_30 <= 1'b1;
              end
              if(_zz_67[31]) begin
                valid_1_31 <= 1'b1;
              end
              if(_zz_68[0]) begin
                dirty_1_0 <= 1'b0;
              end
              if(_zz_68[1]) begin
                dirty_1_1 <= 1'b0;
              end
              if(_zz_68[2]) begin
                dirty_1_2 <= 1'b0;
              end
              if(_zz_68[3]) begin
                dirty_1_3 <= 1'b0;
              end
              if(_zz_68[4]) begin
                dirty_1_4 <= 1'b0;
              end
              if(_zz_68[5]) begin
                dirty_1_5 <= 1'b0;
              end
              if(_zz_68[6]) begin
                dirty_1_6 <= 1'b0;
              end
              if(_zz_68[7]) begin
                dirty_1_7 <= 1'b0;
              end
              if(_zz_68[8]) begin
                dirty_1_8 <= 1'b0;
              end
              if(_zz_68[9]) begin
                dirty_1_9 <= 1'b0;
              end
              if(_zz_68[10]) begin
                dirty_1_10 <= 1'b0;
              end
              if(_zz_68[11]) begin
                dirty_1_11 <= 1'b0;
              end
              if(_zz_68[12]) begin
                dirty_1_12 <= 1'b0;
              end
              if(_zz_68[13]) begin
                dirty_1_13 <= 1'b0;
              end
              if(_zz_68[14]) begin
                dirty_1_14 <= 1'b0;
              end
              if(_zz_68[15]) begin
                dirty_1_15 <= 1'b0;
              end
              if(_zz_68[16]) begin
                dirty_1_16 <= 1'b0;
              end
              if(_zz_68[17]) begin
                dirty_1_17 <= 1'b0;
              end
              if(_zz_68[18]) begin
                dirty_1_18 <= 1'b0;
              end
              if(_zz_68[19]) begin
                dirty_1_19 <= 1'b0;
              end
              if(_zz_68[20]) begin
                dirty_1_20 <= 1'b0;
              end
              if(_zz_68[21]) begin
                dirty_1_21 <= 1'b0;
              end
              if(_zz_68[22]) begin
                dirty_1_22 <= 1'b0;
              end
              if(_zz_68[23]) begin
                dirty_1_23 <= 1'b0;
              end
              if(_zz_68[24]) begin
                dirty_1_24 <= 1'b0;
              end
              if(_zz_68[25]) begin
                dirty_1_25 <= 1'b0;
              end
              if(_zz_68[26]) begin
                dirty_1_26 <= 1'b0;
              end
              if(_zz_68[27]) begin
                dirty_1_27 <= 1'b0;
              end
              if(_zz_68[28]) begin
                dirty_1_28 <= 1'b0;
              end
              if(_zz_68[29]) begin
                dirty_1_29 <= 1'b0;
              end
              if(_zz_68[30]) begin
                dirty_1_30 <= 1'b0;
              end
              if(_zz_68[31]) begin
                dirty_1_31 <= 1'b0;
              end
            end
            if(when_LSU_l473_2) begin
              if(_zz_69[0]) begin
                valid_2_0 <= 1'b1;
              end
              if(_zz_69[1]) begin
                valid_2_1 <= 1'b1;
              end
              if(_zz_69[2]) begin
                valid_2_2 <= 1'b1;
              end
              if(_zz_69[3]) begin
                valid_2_3 <= 1'b1;
              end
              if(_zz_69[4]) begin
                valid_2_4 <= 1'b1;
              end
              if(_zz_69[5]) begin
                valid_2_5 <= 1'b1;
              end
              if(_zz_69[6]) begin
                valid_2_6 <= 1'b1;
              end
              if(_zz_69[7]) begin
                valid_2_7 <= 1'b1;
              end
              if(_zz_69[8]) begin
                valid_2_8 <= 1'b1;
              end
              if(_zz_69[9]) begin
                valid_2_9 <= 1'b1;
              end
              if(_zz_69[10]) begin
                valid_2_10 <= 1'b1;
              end
              if(_zz_69[11]) begin
                valid_2_11 <= 1'b1;
              end
              if(_zz_69[12]) begin
                valid_2_12 <= 1'b1;
              end
              if(_zz_69[13]) begin
                valid_2_13 <= 1'b1;
              end
              if(_zz_69[14]) begin
                valid_2_14 <= 1'b1;
              end
              if(_zz_69[15]) begin
                valid_2_15 <= 1'b1;
              end
              if(_zz_69[16]) begin
                valid_2_16 <= 1'b1;
              end
              if(_zz_69[17]) begin
                valid_2_17 <= 1'b1;
              end
              if(_zz_69[18]) begin
                valid_2_18 <= 1'b1;
              end
              if(_zz_69[19]) begin
                valid_2_19 <= 1'b1;
              end
              if(_zz_69[20]) begin
                valid_2_20 <= 1'b1;
              end
              if(_zz_69[21]) begin
                valid_2_21 <= 1'b1;
              end
              if(_zz_69[22]) begin
                valid_2_22 <= 1'b1;
              end
              if(_zz_69[23]) begin
                valid_2_23 <= 1'b1;
              end
              if(_zz_69[24]) begin
                valid_2_24 <= 1'b1;
              end
              if(_zz_69[25]) begin
                valid_2_25 <= 1'b1;
              end
              if(_zz_69[26]) begin
                valid_2_26 <= 1'b1;
              end
              if(_zz_69[27]) begin
                valid_2_27 <= 1'b1;
              end
              if(_zz_69[28]) begin
                valid_2_28 <= 1'b1;
              end
              if(_zz_69[29]) begin
                valid_2_29 <= 1'b1;
              end
              if(_zz_69[30]) begin
                valid_2_30 <= 1'b1;
              end
              if(_zz_69[31]) begin
                valid_2_31 <= 1'b1;
              end
              if(_zz_70[0]) begin
                dirty_2_0 <= 1'b0;
              end
              if(_zz_70[1]) begin
                dirty_2_1 <= 1'b0;
              end
              if(_zz_70[2]) begin
                dirty_2_2 <= 1'b0;
              end
              if(_zz_70[3]) begin
                dirty_2_3 <= 1'b0;
              end
              if(_zz_70[4]) begin
                dirty_2_4 <= 1'b0;
              end
              if(_zz_70[5]) begin
                dirty_2_5 <= 1'b0;
              end
              if(_zz_70[6]) begin
                dirty_2_6 <= 1'b0;
              end
              if(_zz_70[7]) begin
                dirty_2_7 <= 1'b0;
              end
              if(_zz_70[8]) begin
                dirty_2_8 <= 1'b0;
              end
              if(_zz_70[9]) begin
                dirty_2_9 <= 1'b0;
              end
              if(_zz_70[10]) begin
                dirty_2_10 <= 1'b0;
              end
              if(_zz_70[11]) begin
                dirty_2_11 <= 1'b0;
              end
              if(_zz_70[12]) begin
                dirty_2_12 <= 1'b0;
              end
              if(_zz_70[13]) begin
                dirty_2_13 <= 1'b0;
              end
              if(_zz_70[14]) begin
                dirty_2_14 <= 1'b0;
              end
              if(_zz_70[15]) begin
                dirty_2_15 <= 1'b0;
              end
              if(_zz_70[16]) begin
                dirty_2_16 <= 1'b0;
              end
              if(_zz_70[17]) begin
                dirty_2_17 <= 1'b0;
              end
              if(_zz_70[18]) begin
                dirty_2_18 <= 1'b0;
              end
              if(_zz_70[19]) begin
                dirty_2_19 <= 1'b0;
              end
              if(_zz_70[20]) begin
                dirty_2_20 <= 1'b0;
              end
              if(_zz_70[21]) begin
                dirty_2_21 <= 1'b0;
              end
              if(_zz_70[22]) begin
                dirty_2_22 <= 1'b0;
              end
              if(_zz_70[23]) begin
                dirty_2_23 <= 1'b0;
              end
              if(_zz_70[24]) begin
                dirty_2_24 <= 1'b0;
              end
              if(_zz_70[25]) begin
                dirty_2_25 <= 1'b0;
              end
              if(_zz_70[26]) begin
                dirty_2_26 <= 1'b0;
              end
              if(_zz_70[27]) begin
                dirty_2_27 <= 1'b0;
              end
              if(_zz_70[28]) begin
                dirty_2_28 <= 1'b0;
              end
              if(_zz_70[29]) begin
                dirty_2_29 <= 1'b0;
              end
              if(_zz_70[30]) begin
                dirty_2_30 <= 1'b0;
              end
              if(_zz_70[31]) begin
                dirty_2_31 <= 1'b0;
              end
            end
            if(when_LSU_l473_3) begin
              if(_zz_71[0]) begin
                valid_3_0 <= 1'b1;
              end
              if(_zz_71[1]) begin
                valid_3_1 <= 1'b1;
              end
              if(_zz_71[2]) begin
                valid_3_2 <= 1'b1;
              end
              if(_zz_71[3]) begin
                valid_3_3 <= 1'b1;
              end
              if(_zz_71[4]) begin
                valid_3_4 <= 1'b1;
              end
              if(_zz_71[5]) begin
                valid_3_5 <= 1'b1;
              end
              if(_zz_71[6]) begin
                valid_3_6 <= 1'b1;
              end
              if(_zz_71[7]) begin
                valid_3_7 <= 1'b1;
              end
              if(_zz_71[8]) begin
                valid_3_8 <= 1'b1;
              end
              if(_zz_71[9]) begin
                valid_3_9 <= 1'b1;
              end
              if(_zz_71[10]) begin
                valid_3_10 <= 1'b1;
              end
              if(_zz_71[11]) begin
                valid_3_11 <= 1'b1;
              end
              if(_zz_71[12]) begin
                valid_3_12 <= 1'b1;
              end
              if(_zz_71[13]) begin
                valid_3_13 <= 1'b1;
              end
              if(_zz_71[14]) begin
                valid_3_14 <= 1'b1;
              end
              if(_zz_71[15]) begin
                valid_3_15 <= 1'b1;
              end
              if(_zz_71[16]) begin
                valid_3_16 <= 1'b1;
              end
              if(_zz_71[17]) begin
                valid_3_17 <= 1'b1;
              end
              if(_zz_71[18]) begin
                valid_3_18 <= 1'b1;
              end
              if(_zz_71[19]) begin
                valid_3_19 <= 1'b1;
              end
              if(_zz_71[20]) begin
                valid_3_20 <= 1'b1;
              end
              if(_zz_71[21]) begin
                valid_3_21 <= 1'b1;
              end
              if(_zz_71[22]) begin
                valid_3_22 <= 1'b1;
              end
              if(_zz_71[23]) begin
                valid_3_23 <= 1'b1;
              end
              if(_zz_71[24]) begin
                valid_3_24 <= 1'b1;
              end
              if(_zz_71[25]) begin
                valid_3_25 <= 1'b1;
              end
              if(_zz_71[26]) begin
                valid_3_26 <= 1'b1;
              end
              if(_zz_71[27]) begin
                valid_3_27 <= 1'b1;
              end
              if(_zz_71[28]) begin
                valid_3_28 <= 1'b1;
              end
              if(_zz_71[29]) begin
                valid_3_29 <= 1'b1;
              end
              if(_zz_71[30]) begin
                valid_3_30 <= 1'b1;
              end
              if(_zz_71[31]) begin
                valid_3_31 <= 1'b1;
              end
              if(_zz_72[0]) begin
                dirty_3_0 <= 1'b0;
              end
              if(_zz_72[1]) begin
                dirty_3_1 <= 1'b0;
              end
              if(_zz_72[2]) begin
                dirty_3_2 <= 1'b0;
              end
              if(_zz_72[3]) begin
                dirty_3_3 <= 1'b0;
              end
              if(_zz_72[4]) begin
                dirty_3_4 <= 1'b0;
              end
              if(_zz_72[5]) begin
                dirty_3_5 <= 1'b0;
              end
              if(_zz_72[6]) begin
                dirty_3_6 <= 1'b0;
              end
              if(_zz_72[7]) begin
                dirty_3_7 <= 1'b0;
              end
              if(_zz_72[8]) begin
                dirty_3_8 <= 1'b0;
              end
              if(_zz_72[9]) begin
                dirty_3_9 <= 1'b0;
              end
              if(_zz_72[10]) begin
                dirty_3_10 <= 1'b0;
              end
              if(_zz_72[11]) begin
                dirty_3_11 <= 1'b0;
              end
              if(_zz_72[12]) begin
                dirty_3_12 <= 1'b0;
              end
              if(_zz_72[13]) begin
                dirty_3_13 <= 1'b0;
              end
              if(_zz_72[14]) begin
                dirty_3_14 <= 1'b0;
              end
              if(_zz_72[15]) begin
                dirty_3_15 <= 1'b0;
              end
              if(_zz_72[16]) begin
                dirty_3_16 <= 1'b0;
              end
              if(_zz_72[17]) begin
                dirty_3_17 <= 1'b0;
              end
              if(_zz_72[18]) begin
                dirty_3_18 <= 1'b0;
              end
              if(_zz_72[19]) begin
                dirty_3_19 <= 1'b0;
              end
              if(_zz_72[20]) begin
                dirty_3_20 <= 1'b0;
              end
              if(_zz_72[21]) begin
                dirty_3_21 <= 1'b0;
              end
              if(_zz_72[22]) begin
                dirty_3_22 <= 1'b0;
              end
              if(_zz_72[23]) begin
                dirty_3_23 <= 1'b0;
              end
              if(_zz_72[24]) begin
                dirty_3_24 <= 1'b0;
              end
              if(_zz_72[25]) begin
                dirty_3_25 <= 1'b0;
              end
              if(_zz_72[26]) begin
                dirty_3_26 <= 1'b0;
              end
              if(_zz_72[27]) begin
                dirty_3_27 <= 1'b0;
              end
              if(_zz_72[28]) begin
                dirty_3_28 <= 1'b0;
              end
              if(_zz_72[29]) begin
                dirty_3_29 <= 1'b0;
              end
              if(_zz_72[30]) begin
                dirty_3_30 <= 1'b0;
              end
              if(_zz_72[31]) begin
                dirty_3_31 <= 1'b0;
              end
            end
          end
        end
        axiCtrl_enumDef_readFirst : begin
          if(when_LSU_l496) begin
            transferRAddrMid <= _zz_transferRAddrMid;
          end
        end
        axiCtrl_enumDef_read : begin
          if(when_LSU_l510) begin
            transferRAddrMid <= _zz_transferRAddrMid_1;
          end
        end
        axiCtrl_enumDef_writeReq : begin
        end
        axiCtrl_enumDef_write : begin
          if(when_LSU_l539) begin
            transferWAddrMid <= _zz_transferWAddrMid;
            if(io_axi_wlast) begin
              if(!transferUncached) begin
                if(transferCACOP) begin
                  transferCACOP <= 1'b0;
                end
              end
            end
          end
        end
        default : begin
        end
      endcase
      rollbackCtrl_stateReg <= rollbackCtrl_stateNext;
      case(rollbackCtrl_stateReg)
        rollbackCtrl_enumDef_idle : begin
          if(when_LSU_l564) begin
            writeBufferTail <= (writeBufferTail + 3'b001);
          end
          if(when_LSU_l567) begin
            writeBufferTail <= (writeBufferTail - 3'b001);
          end
        end
        rollbackCtrl_enumDef_rollback : begin
          if(!when_LSU_l575) begin
            writeBufferTail <= (writeBufferTail - 3'b001);
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge aclk) begin
    if(stage1Out_thrown_ready) begin
      stage1Out_thrown_rData_robIdx <= stage1Out_thrown_payload_robIdx;
      stage1Out_thrown_rData_prd <= stage1Out_thrown_payload_prd;
      stage1Out_thrown_rData_branchResult_targetPC <= stage1Out_thrown_payload_branchResult_targetPC;
      stage1Out_thrown_rData_branchResult_branchResult <= stage1Out_thrown_payload_branchResult_branchResult;
      stage1Out_thrown_rData_branchResult_predictFail <= stage1Out_thrown_payload_branchResult_predictFail;
      stage1Out_thrown_rData_exceptionInfo_exception <= stage1Out_thrown_payload_exceptionInfo_exception;
      stage1Out_thrown_rData_exceptionInfo_eCode <= stage1Out_thrown_payload_exceptionInfo_eCode;
      stage1Out_thrown_rData_exceptionInfo_eSubCode <= stage1Out_thrown_payload_exceptionInfo_eSubCode;
      stage1Out_thrown_rData_storeData <= stage1Out_thrown_payload_storeData;
      stage1Out_thrown_rData_lsCtrlBundle_load <= stage1Out_thrown_payload_lsCtrlBundle_load;
      stage1Out_thrown_rData_lsCtrlBundle_store <= stage1Out_thrown_payload_lsCtrlBundle_store;
      stage1Out_thrown_rData_lsCtrlBundle_signed <= stage1Out_thrown_payload_lsCtrlBundle_signed;
      stage1Out_thrown_rData_lsCtrlBundle_ll <= stage1Out_thrown_payload_lsCtrlBundle_ll;
      stage1Out_thrown_rData_lsCtrlBundle_sc <= stage1Out_thrown_payload_lsCtrlBundle_sc;
      stage1Out_thrown_rData_lsCtrlBundle_lsMask <= stage1Out_thrown_payload_lsCtrlBundle_lsMask;
      stage1Out_thrown_rData_lsCtrlBundle_size <= stage1Out_thrown_payload_lsCtrlBundle_size;
      stage1Out_thrown_rData_lsCtrlBundle_normalMemOp <= stage1Out_thrown_payload_lsCtrlBundle_normalMemOp;
      stage1Out_thrown_rData_vaddr <= stage1Out_thrown_payload_vaddr;
      stage1Out_thrown_rData_tlb_hit <= stage1Out_thrown_payload_tlb_hit;
      stage1Out_thrown_rData_tlb_pageInfo_ppn <= stage1Out_thrown_payload_tlb_pageInfo_ppn;
      stage1Out_thrown_rData_tlb_pageInfo_plv <= stage1Out_thrown_payload_tlb_pageInfo_plv;
      stage1Out_thrown_rData_tlb_pageInfo_mat <= stage1Out_thrown_payload_tlb_pageInfo_mat;
      stage1Out_thrown_rData_tlb_pageInfo_d <= stage1Out_thrown_payload_tlb_pageInfo_d;
      stage1Out_thrown_rData_tlb_pageInfo_v <= stage1Out_thrown_payload_tlb_pageInfo_v;
      stage1Out_thrown_rData_wayValid <= stage1Out_thrown_payload_wayValid;
      stage1Out_thrown_rData_wayDirty <= stage1Out_thrown_payload_wayDirty;
      stage1Out_thrown_rData_isStoreTag <= stage1Out_thrown_payload_isStoreTag;
      stage1Out_thrown_rData_isIndexInvalidate <= stage1Out_thrown_payload_isIndexInvalidate;
      stage1Out_thrown_rData_isHitInvalidate <= stage1Out_thrown_payload_isHitInvalidate;
      stage1Out_thrown_rData_checkTLBException <= stage1Out_thrown_payload_checkTLBException;
      stage1Out_thrown_rData_lsException <= stage1Out_thrown_payload_lsException;
    end
  end


endmodule

module ICache (
  input  wire          io_input_0_valid,
  output wire          io_input_0_ready,
  input  wire [31:0]   io_input_0_payload_address,
  input  wire [3:0]    io_input_0_payload_size,
  input  wire [31:0]   io_input_0_payload_branchInfo_predictPC,
  input  wire          io_input_0_payload_branchInfo_predictResult,
  input  wire          io_input_1_valid,
  output wire          io_input_1_ready,
  input  wire [31:0]   io_input_1_payload_address,
  input  wire [3:0]    io_input_1_payload_size,
  input  wire [31:0]   io_input_1_payload_branchInfo_predictPC,
  input  wire          io_input_1_payload_branchInfo_predictResult,
  input  wire [1:0]    io_output_allowMask,
  output wire [1:0]    io_output_availMask,
  output wire [31:0]   io_output_info_0_inst,
  output wire [31:0]   io_output_info_0_branchInfo_predictPC,
  output wire          io_output_info_0_branchInfo_predictResult,
  output wire          io_output_info_0_exceptionInfo_exception,
  output wire [5:0]    io_output_info_0_exceptionInfo_eCode,
  output wire [0:0]    io_output_info_0_exceptionInfo_eSubCode,
  output wire [31:0]   io_output_info_0_pc,
  output wire [31:0]   io_output_info_1_inst,
  output wire [31:0]   io_output_info_1_branchInfo_predictPC,
  output wire          io_output_info_1_branchInfo_predictResult,
  output wire          io_output_info_1_exceptionInfo_exception,
  output wire [5:0]    io_output_info_1_exceptionInfo_eCode,
  output wire [0:0]    io_output_info_1_exceptionInfo_eSubCode,
  output wire [31:0]   io_output_info_1_pc,
  input  wire          io_tlb_hit,
  input  wire [19:0]   io_tlb_pageInfo_ppn,
  input  wire [1:0]    io_tlb_pageInfo_plv,
  input  wire [1:0]    io_tlb_pageInfo_mat,
  input  wire          io_tlb_pageInfo_d,
  input  wire          io_tlb_pageInfo_v,
  output wire [19:0]   io_tlb_virtPageNumber,
  input  wire [1:0]    _zz_when_Cache_l83,
  output wire          io_ctrl_busy,
  input  wire          io_ctrl_stall,
  input  wire [31:0]   io_ctrl_cacopVA,
  input  wire          io_ctrl_cacopStoreTag,
  input  wire          io_ctrl_cacopIndexInvalidate,
  input  wire          io_ctrl_cacopHitInvalidate,
  input  wire          io_flush,
  output wire [31:0]   io_badv_vaddr,
  output wire          io_badv_wen,
  output wire [3:0]    io_axi_arid,
  output wire [31:0]   io_axi_araddr,
  output wire [7:0]    io_axi_arlen,
  output wire [2:0]    io_axi_arsize,
  output wire [1:0]    io_axi_arburst,
  output wire [1:0]    io_axi_arlock,
  output wire [3:0]    io_axi_arcache,
  output wire [2:0]    io_axi_arprot,
  output reg           io_axi_arvalid,
  input  wire          io_axi_arready,
  input  wire [3:0]    io_axi_rid,
  input  wire [31:0]   io_axi_rdata,
  input  wire [1:0]    io_axi_rresp,
  input  wire          io_axi_rlast,
  input  wire          io_axi_rvalid,
  output reg           io_axi_rready,
  input  wire          aclk,
  input  wire          aresetn
);
  localparam LSUSizeOp_byte_1 = 4'd1;
  localparam LSUSizeOp_halfword = 4'd3;
  localparam LSUSizeOp_word = 4'd15;
  localparam fsm_enumDef_1_BOOT = 2'd0;
  localparam fsm_enumDef_1_idle = 2'd1;
  localparam fsm_enumDef_1_req = 2'd2;
  localparam fsm_enumDef_1_read = 2'd3;

  wire                data_0_wr_en;
  wire       [0:0]    data_0_wr_mask;
  wire                data_0_rd_en;
  wire       [8:0]    data_0_rd_addr;
  wire                data_0_1_wr_en;
  wire       [0:0]    data_0_1_wr_mask;
  wire                data_0_1_rd_en;
  wire       [8:0]    data_0_1_rd_addr;
  wire                data_1_wr_en;
  wire       [0:0]    data_1_wr_mask;
  wire                data_1_rd_en;
  wire       [8:0]    data_1_rd_addr;
  wire                data_1_1_wr_en;
  wire       [0:0]    data_1_1_wr_mask;
  wire                data_1_1_rd_en;
  wire       [8:0]    data_1_1_rd_addr;
  wire                data_2_wr_en;
  wire       [0:0]    data_2_wr_mask;
  wire                data_2_rd_en;
  wire       [8:0]    data_2_rd_addr;
  wire                data_2_1_wr_en;
  wire       [0:0]    data_2_1_wr_mask;
  wire                data_2_1_rd_en;
  wire       [8:0]    data_2_1_rd_addr;
  wire                data_3_wr_en;
  wire       [0:0]    data_3_wr_mask;
  wire                data_3_rd_en;
  wire       [8:0]    data_3_rd_addr;
  wire                data_3_1_wr_en;
  wire       [0:0]    data_3_1_wr_mask;
  wire                data_3_1_rd_en;
  wire       [8:0]    data_3_1_rd_addr;
  wire                tag_0_wr_en;
  wire       [0:0]    tag_0_wr_mask;
  wire                tag_0_rd_en;
  wire       [4:0]    tag_0_rd_addr;
  wire                tag_0_1_wr_en;
  wire       [0:0]    tag_0_1_wr_mask;
  wire                tag_0_1_rd_en;
  wire       [4:0]    tag_0_1_rd_addr;
  wire                tag_1_wr_en;
  wire       [0:0]    tag_1_wr_mask;
  wire                tag_1_rd_en;
  wire       [4:0]    tag_1_rd_addr;
  wire                tag_1_1_wr_en;
  wire       [0:0]    tag_1_1_wr_mask;
  wire                tag_1_1_rd_en;
  wire       [4:0]    tag_1_1_rd_addr;
  wire                tag_2_wr_en;
  wire       [0:0]    tag_2_wr_mask;
  wire                tag_2_rd_en;
  wire       [4:0]    tag_2_rd_addr;
  wire                tag_2_1_wr_en;
  wire       [0:0]    tag_2_1_wr_mask;
  wire                tag_2_1_rd_en;
  wire       [4:0]    tag_2_1_rd_addr;
  wire                tag_3_wr_en;
  wire       [0:0]    tag_3_wr_mask;
  wire                tag_3_rd_en;
  wire       [4:0]    tag_3_rd_addr;
  wire                tag_3_1_wr_en;
  wire       [0:0]    tag_3_1_wr_mask;
  wire                tag_3_1_rd_en;
  wire       [4:0]    tag_3_1_rd_addr;
  wire       [31:0]   data_0_rd_data;
  wire       [31:0]   data_0_1_rd_data;
  wire       [31:0]   data_1_rd_data;
  wire       [31:0]   data_1_1_rd_data;
  wire       [31:0]   data_2_rd_data;
  wire       [31:0]   data_2_1_rd_data;
  wire       [31:0]   data_3_rd_data;
  wire       [31:0]   data_3_1_rd_data;
  wire       [20:0]   tag_0_rd_data;
  wire       [20:0]   tag_0_1_rd_data;
  wire       [20:0]   tag_1_rd_data;
  wire       [20:0]   tag_1_1_rd_data;
  wire       [20:0]   tag_2_rd_data;
  wire       [20:0]   tag_2_1_rd_data;
  wire       [20:0]   tag_3_rd_data;
  wire       [20:0]   tag_3_1_rd_data;
  wire       [1:0]    _zz_acceptMask;
  reg        [1:0]    _zz_acceptMask_1;
  wire       [1:0]    _zz_acceptMask_2;
  reg                 _zz_stage1Out_payload_wayValid_0;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_0_1;
  wire       [31:0]   _zz_stage1Out_payload_wayValid_0_2;
  wire       [1:0]    _zz_hit_0;
  wire       [0:0]    _zz_hit_0_1;
  reg                 _zz_stage1Out_payload_wayValid_0_3;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_0_4;
  wire       [31:0]   _zz_stage1Out_payload_wayValid_0_5;
  wire       [1:0]    _zz_hit_0_2;
  wire       [0:0]    _zz_hit_0_3;
  reg                 _zz_stage1Out_payload_wayValid_0_6;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_0_7;
  wire       [31:0]   _zz_stage1Out_payload_wayValid_0_8;
  wire       [1:0]    _zz_hit_0_4;
  wire       [0:0]    _zz_hit_0_5;
  reg                 _zz_stage1Out_payload_wayValid_0_9;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_0_10;
  wire       [31:0]   _zz_stage1Out_payload_wayValid_0_11;
  wire       [1:0]    _zz_hit_0_6;
  wire       [0:0]    _zz_hit_0_7;
  reg                 _zz_stage1Out_payload_wayValid_1;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_1_1;
  wire       [1:0]    _zz_hit_1;
  wire       [0:0]    _zz_hit_1_1;
  reg                 _zz_stage1Out_payload_wayValid_1_2;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_1_3;
  wire       [1:0]    _zz_hit_1_2;
  wire       [0:0]    _zz_hit_1_3;
  reg                 _zz_stage1Out_payload_wayValid_1_4;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_1_5;
  wire       [1:0]    _zz_hit_1_4;
  wire       [0:0]    _zz_hit_1_5;
  reg                 _zz_stage1Out_payload_wayValid_1_6;
  wire       [4:0]    _zz_stage1Out_payload_wayValid_1_7;
  wire       [1:0]    _zz_hit_1_6;
  wire       [0:0]    _zz_hit_1_7;
  reg        [1:0]    _zz_fireMask;
  wire       [1:0]    _zz_fireMask_1;
  wire       [1:0]    _zz_exceptionInfo2_eCode;
  wire       [2:0]    _zz_exceptionInfo2_eCode_1;
  wire       [2:0]    _zz_exceptionInfo2_eCode_2;
  wire       [1:0]    _zz_when_Cache_l131;
  wire       [0:0]    _zz_when_Cache_l131_1;
  wire       [1:0]    _zz_when_Cache_l131_1_1;
  wire       [0:0]    _zz_when_Cache_l131_1_2;
  wire       [7:0]    _zz_io_axi_arlen;
  wire       [3:0]    _zz_io_axi_arlen_1;
  wire       [3:0]    _zz_exceptionInfo1_0_eCode;
  wire       [3:0]    _zz_exceptionInfo1_0_eCode_1;
  reg        [31:0]   _zz_portData_0_inst_3;
  wire       [1:0]    _zz_portData_0_inst_4;
  wire       [1:0]    _zz__zz_io_output_info_0_inst;
  reg        [1:0]    _zz__zz_io_output_info_0_inst_1;
  wire       [1:0]    _zz__zz_io_output_info_0_inst_2;
  reg        [31:0]   _zz_io_output_info_0_inst_1;
  reg        [31:0]   _zz_io_output_info_0_branchInfo_predictPC;
  reg                 _zz_io_output_info_0_branchInfo_predictResult;
  reg                 _zz_io_output_info_0_exceptionInfo_exception;
  reg        [5:0]    _zz_io_output_info_0_exceptionInfo_eCode;
  reg        [0:0]    _zz_io_output_info_0_exceptionInfo_eSubCode;
  reg        [31:0]   _zz_io_output_info_0_pc;
  reg                 _zz__zz_wayToReplace_0;
  wire       [4:0]    _zz__zz_wayToReplace_0_1;
  reg                 _zz__zz_wayToReplace_0_2;
  wire       [4:0]    _zz__zz_wayToReplace_0_3;
  reg                 _zz__zz_wayToReplace_0_1_1;
  wire       [4:0]    _zz__zz_wayToReplace_0_1_2;
  reg                 _zz__zz_wayToReplace_0_1_3;
  wire       [4:0]    _zz__zz_wayToReplace_0_1_4;
  reg                 _zz__zz_wayToReplace_0_2_1;
  wire       [4:0]    _zz__zz_wayToReplace_0_2_2;
  reg                 _zz__zz_wayToReplace_0_2_3;
  wire       [4:0]    _zz__zz_wayToReplace_0_2_4;
  reg                 _zz__zz_wayToReplace_0_3_1;
  wire       [4:0]    _zz__zz_wayToReplace_0_3_2;
  reg                 _zz__zz_wayToReplace_0_3_3;
  wire       [4:0]    _zz__zz_wayToReplace_0_3_4;
  wire       [3:0]    _zz_exceptionInfo1_1_eCode;
  wire       [3:0]    _zz_exceptionInfo1_1_eCode_1;
  reg        [31:0]   _zz_portData_1_inst_3;
  wire       [1:0]    _zz_portData_1_inst_4;
  wire       [1:0]    _zz__zz_io_output_info_1_inst;
  reg        [1:0]    _zz__zz_io_output_info_1_inst_1;
  wire       [1:0]    _zz__zz_io_output_info_1_inst_2;
  reg        [31:0]   _zz_io_output_info_1_inst_1;
  reg        [31:0]   _zz_io_output_info_1_branchInfo_predictPC;
  reg                 _zz_io_output_info_1_branchInfo_predictResult;
  reg                 _zz_io_output_info_1_exceptionInfo_exception;
  reg        [5:0]    _zz_io_output_info_1_exceptionInfo_eCode;
  reg        [0:0]    _zz_io_output_info_1_exceptionInfo_eSubCode;
  reg        [31:0]   _zz_io_output_info_1_pc;
  reg                 _zz__zz_wayToReplace_1;
  wire       [4:0]    _zz__zz_wayToReplace_1_1;
  reg                 _zz__zz_wayToReplace_1_2;
  wire       [4:0]    _zz__zz_wayToReplace_1_3;
  reg                 _zz__zz_wayToReplace_1_1_1;
  wire       [4:0]    _zz__zz_wayToReplace_1_1_2;
  reg                 _zz__zz_wayToReplace_1_1_3;
  wire       [4:0]    _zz__zz_wayToReplace_1_1_4;
  reg                 _zz__zz_wayToReplace_1_2_1;
  wire       [4:0]    _zz__zz_wayToReplace_1_2_2;
  reg                 _zz__zz_wayToReplace_1_2_3;
  wire       [4:0]    _zz__zz_wayToReplace_1_2_4;
  reg                 _zz__zz_wayToReplace_1_3_1;
  wire       [4:0]    _zz__zz_wayToReplace_1_3_2;
  reg                 _zz__zz_wayToReplace_1_3_3;
  wire       [4:0]    _zz__zz_wayToReplace_1_3_4;
  reg        [1:0]    _zz_io_output_availMask_2;
  wire       [1:0]    _zz_io_output_availMask_3;
  wire       [3:0]    _zz_cacopWay;
  wire       [1:0]    _zz_when_Cache_l198;
  wire       [0:0]    _zz_when_Cache_l198_1;
  wire       [1:0]    _zz_when_Cache_l180;
  wire       [0:0]    _zz_when_Cache_l180_1;
  wire       [31:0]   _zz_rd_addr;
  wire       [31:0]   _zz_rd_addr_1;
  wire       [31:0]   _zz_rd_addr_2;
  wire       [31:0]   _zz_rd_addr_3;
  wire       [31:0]   _zz_rd_addr_4;
  wire       [31:0]   _zz_rd_addr_5;
  wire       [31:0]   _zz_rd_addr_6;
  wire       [31:0]   _zz_rd_addr_7;
  reg                 _zz_wr_en;
  reg                 _zz_wr_en_1;
  reg                 _zz_wr_en_2;
  reg                 _zz_wr_en_3;
  reg                 _zz_wr_en_4;
  reg                 _zz_wr_en_5;
  reg                 _zz_wr_en_6;
  reg                 _zz_wr_en_7;
  reg                 valid_0_0;
  reg                 valid_0_1;
  reg                 valid_0_2;
  reg                 valid_0_3;
  reg                 valid_0_4;
  reg                 valid_0_5;
  reg                 valid_0_6;
  reg                 valid_0_7;
  reg                 valid_0_8;
  reg                 valid_0_9;
  reg                 valid_0_10;
  reg                 valid_0_11;
  reg                 valid_0_12;
  reg                 valid_0_13;
  reg                 valid_0_14;
  reg                 valid_0_15;
  reg                 valid_0_16;
  reg                 valid_0_17;
  reg                 valid_0_18;
  reg                 valid_0_19;
  reg                 valid_0_20;
  reg                 valid_0_21;
  reg                 valid_0_22;
  reg                 valid_0_23;
  reg                 valid_0_24;
  reg                 valid_0_25;
  reg                 valid_0_26;
  reg                 valid_0_27;
  reg                 valid_0_28;
  reg                 valid_0_29;
  reg                 valid_0_30;
  reg                 valid_0_31;
  reg                 valid_1_0;
  reg                 valid_1_1;
  reg                 valid_1_2;
  reg                 valid_1_3;
  reg                 valid_1_4;
  reg                 valid_1_5;
  reg                 valid_1_6;
  reg                 valid_1_7;
  reg                 valid_1_8;
  reg                 valid_1_9;
  reg                 valid_1_10;
  reg                 valid_1_11;
  reg                 valid_1_12;
  reg                 valid_1_13;
  reg                 valid_1_14;
  reg                 valid_1_15;
  reg                 valid_1_16;
  reg                 valid_1_17;
  reg                 valid_1_18;
  reg                 valid_1_19;
  reg                 valid_1_20;
  reg                 valid_1_21;
  reg                 valid_1_22;
  reg                 valid_1_23;
  reg                 valid_1_24;
  reg                 valid_1_25;
  reg                 valid_1_26;
  reg                 valid_1_27;
  reg                 valid_1_28;
  reg                 valid_1_29;
  reg                 valid_1_30;
  reg                 valid_1_31;
  reg                 valid_2_0;
  reg                 valid_2_1;
  reg                 valid_2_2;
  reg                 valid_2_3;
  reg                 valid_2_4;
  reg                 valid_2_5;
  reg                 valid_2_6;
  reg                 valid_2_7;
  reg                 valid_2_8;
  reg                 valid_2_9;
  reg                 valid_2_10;
  reg                 valid_2_11;
  reg                 valid_2_12;
  reg                 valid_2_13;
  reg                 valid_2_14;
  reg                 valid_2_15;
  reg                 valid_2_16;
  reg                 valid_2_17;
  reg                 valid_2_18;
  reg                 valid_2_19;
  reg                 valid_2_20;
  reg                 valid_2_21;
  reg                 valid_2_22;
  reg                 valid_2_23;
  reg                 valid_2_24;
  reg                 valid_2_25;
  reg                 valid_2_26;
  reg                 valid_2_27;
  reg                 valid_2_28;
  reg                 valid_2_29;
  reg                 valid_2_30;
  reg                 valid_2_31;
  reg                 valid_3_0;
  reg                 valid_3_1;
  reg                 valid_3_2;
  reg                 valid_3_3;
  reg                 valid_3_4;
  reg                 valid_3_5;
  reg                 valid_3_6;
  reg                 valid_3_7;
  reg                 valid_3_8;
  reg                 valid_3_9;
  reg                 valid_3_10;
  reg                 valid_3_11;
  reg                 valid_3_12;
  reg                 valid_3_13;
  reg                 valid_3_14;
  reg                 valid_3_15;
  reg                 valid_3_16;
  reg                 valid_3_17;
  reg                 valid_3_18;
  reg                 valid_3_19;
  reg                 valid_3_20;
  reg                 valid_3_21;
  reg                 valid_3_22;
  reg                 valid_3_23;
  reg                 valid_3_24;
  reg                 valid_3_25;
  reg                 valid_3_26;
  reg                 valid_3_27;
  reg                 valid_3_28;
  reg                 valid_3_29;
  reg                 valid_3_30;
  reg                 valid_3_31;
  wire       [31:0]   dataRead_0_0;
  wire       [31:0]   dataRead_0_1;
  wire       [31:0]   dataRead_0_2;
  wire       [31:0]   dataRead_0_3;
  wire       [31:0]   dataRead_1_0;
  wire       [31:0]   dataRead_1_1;
  wire       [31:0]   dataRead_1_2;
  wire       [31:0]   dataRead_1_3;
  wire       [20:0]   tagRead_0_0;
  wire       [20:0]   tagRead_0_1;
  wire       [20:0]   tagRead_0_2;
  wire       [20:0]   tagRead_0_3;
  wire       [20:0]   tagRead_1_0;
  wire       [20:0]   tagRead_1_1;
  wire       [20:0]   tagRead_1_2;
  wire       [20:0]   tagRead_1_3;
  reg        [3:0]    hit_0;
  reg        [3:0]    hit_1;
  reg        [1:0]    miss;
  wire                stall;
  wire                cacopEn;
  wire                stage1Out_valid;
  reg                 stage1Out_ready;
  wire       [31:0]   stage1Out_payload_branchInfo_0_predictPC;
  wire                stage1Out_payload_branchInfo_0_predictResult;
  wire       [31:0]   stage1Out_payload_branchInfo_1_predictPC;
  wire                stage1Out_payload_branchInfo_1_predictResult;
  wire                stage1Out_payload_exceptionInfo_0_exception;
  wire       [5:0]    stage1Out_payload_exceptionInfo_0_eCode;
  wire       [0:0]    stage1Out_payload_exceptionInfo_0_eSubCode;
  wire                stage1Out_payload_exceptionInfo_1_exception;
  wire       [5:0]    stage1Out_payload_exceptionInfo_1_eCode;
  wire       [0:0]    stage1Out_payload_exceptionInfo_1_eSubCode;
  wire       [31:0]   stage1Out_payload_pc_0;
  wire       [31:0]   stage1Out_payload_pc_1;
  reg        [1:0]    stage1Out_payload_valid;
  wire                stage1Out_payload_tlb_hit;
  wire       [19:0]   stage1Out_payload_tlb_pageInfo_ppn;
  wire       [1:0]    stage1Out_payload_tlb_pageInfo_plv;
  wire       [1:0]    stage1Out_payload_tlb_pageInfo_mat;
  wire                stage1Out_payload_tlb_pageInfo_d;
  wire                stage1Out_payload_tlb_pageInfo_v;
  reg        [3:0]    stage1Out_payload_wayValid_0;
  reg        [3:0]    stage1Out_payload_wayValid_1;
  wire                stage1Out_payload_isStoreTag;
  wire                stage1Out_payload_isIndexInvalidate;
  wire                stage1Out_payload_isHitInvalidate;
  wire                stage2In_valid;
  wire                stage2In_ready;
  wire       [31:0]   stage2In_payload_branchInfo_0_predictPC;
  wire                stage2In_payload_branchInfo_0_predictResult;
  wire       [31:0]   stage2In_payload_branchInfo_1_predictPC;
  wire                stage2In_payload_branchInfo_1_predictResult;
  wire                stage2In_payload_exceptionInfo_0_exception;
  wire       [5:0]    stage2In_payload_exceptionInfo_0_eCode;
  wire       [0:0]    stage2In_payload_exceptionInfo_0_eSubCode;
  wire                stage2In_payload_exceptionInfo_1_exception;
  wire       [5:0]    stage2In_payload_exceptionInfo_1_eCode;
  wire       [0:0]    stage2In_payload_exceptionInfo_1_eSubCode;
  wire       [31:0]   stage2In_payload_pc_0;
  wire       [31:0]   stage2In_payload_pc_1;
  wire       [1:0]    stage2In_payload_valid;
  wire                stage2In_payload_tlb_hit;
  wire       [19:0]   stage2In_payload_tlb_pageInfo_ppn;
  wire       [1:0]    stage2In_payload_tlb_pageInfo_plv;
  wire       [1:0]    stage2In_payload_tlb_pageInfo_mat;
  wire                stage2In_payload_tlb_pageInfo_d;
  wire                stage2In_payload_tlb_pageInfo_v;
  wire       [3:0]    stage2In_payload_wayValid_0;
  wire       [3:0]    stage2In_payload_wayValid_1;
  wire                stage2In_payload_isStoreTag;
  wire                stage2In_payload_isIndexInvalidate;
  wire                stage2In_payload_isHitInvalidate;
  reg                 stage1Out_thrown_valid;
  reg                 stage1Out_thrown_ready;
  wire       [31:0]   stage1Out_thrown_payload_branchInfo_0_predictPC;
  wire                stage1Out_thrown_payload_branchInfo_0_predictResult;
  wire       [31:0]   stage1Out_thrown_payload_branchInfo_1_predictPC;
  wire                stage1Out_thrown_payload_branchInfo_1_predictResult;
  wire                stage1Out_thrown_payload_exceptionInfo_0_exception;
  wire       [5:0]    stage1Out_thrown_payload_exceptionInfo_0_eCode;
  wire       [0:0]    stage1Out_thrown_payload_exceptionInfo_0_eSubCode;
  wire                stage1Out_thrown_payload_exceptionInfo_1_exception;
  wire       [5:0]    stage1Out_thrown_payload_exceptionInfo_1_eCode;
  wire       [0:0]    stage1Out_thrown_payload_exceptionInfo_1_eSubCode;
  wire       [31:0]   stage1Out_thrown_payload_pc_0;
  wire       [31:0]   stage1Out_thrown_payload_pc_1;
  wire       [1:0]    stage1Out_thrown_payload_valid;
  wire                stage1Out_thrown_payload_tlb_hit;
  wire       [19:0]   stage1Out_thrown_payload_tlb_pageInfo_ppn;
  wire       [1:0]    stage1Out_thrown_payload_tlb_pageInfo_plv;
  wire       [1:0]    stage1Out_thrown_payload_tlb_pageInfo_mat;
  wire                stage1Out_thrown_payload_tlb_pageInfo_d;
  wire                stage1Out_thrown_payload_tlb_pageInfo_v;
  wire       [3:0]    stage1Out_thrown_payload_wayValid_0;
  wire       [3:0]    stage1Out_thrown_payload_wayValid_1;
  wire                stage1Out_thrown_payload_isStoreTag;
  wire                stage1Out_thrown_payload_isIndexInvalidate;
  wire                stage1Out_thrown_payload_isHitInvalidate;
  wire                stage1Out_thrown_m2sPipe_valid;
  wire                stage1Out_thrown_m2sPipe_ready;
  wire       [31:0]   stage1Out_thrown_m2sPipe_payload_branchInfo_0_predictPC;
  wire                stage1Out_thrown_m2sPipe_payload_branchInfo_0_predictResult;
  wire       [31:0]   stage1Out_thrown_m2sPipe_payload_branchInfo_1_predictPC;
  wire                stage1Out_thrown_m2sPipe_payload_branchInfo_1_predictResult;
  wire                stage1Out_thrown_m2sPipe_payload_exceptionInfo_0_exception;
  wire       [5:0]    stage1Out_thrown_m2sPipe_payload_exceptionInfo_0_eCode;
  wire       [0:0]    stage1Out_thrown_m2sPipe_payload_exceptionInfo_0_eSubCode;
  wire                stage1Out_thrown_m2sPipe_payload_exceptionInfo_1_exception;
  wire       [5:0]    stage1Out_thrown_m2sPipe_payload_exceptionInfo_1_eCode;
  wire       [0:0]    stage1Out_thrown_m2sPipe_payload_exceptionInfo_1_eSubCode;
  wire       [31:0]   stage1Out_thrown_m2sPipe_payload_pc_0;
  wire       [31:0]   stage1Out_thrown_m2sPipe_payload_pc_1;
  wire       [1:0]    stage1Out_thrown_m2sPipe_payload_valid;
  wire                stage1Out_thrown_m2sPipe_payload_tlb_hit;
  wire       [19:0]   stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_ppn;
  wire       [1:0]    stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_plv;
  wire       [1:0]    stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_mat;
  wire                stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_d;
  wire                stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_v;
  wire       [3:0]    stage1Out_thrown_m2sPipe_payload_wayValid_0;
  wire       [3:0]    stage1Out_thrown_m2sPipe_payload_wayValid_1;
  wire                stage1Out_thrown_m2sPipe_payload_isStoreTag;
  wire                stage1Out_thrown_m2sPipe_payload_isIndexInvalidate;
  wire                stage1Out_thrown_m2sPipe_payload_isHitInvalidate;
  reg                 stage1Out_thrown_rValid;
  reg        [31:0]   stage1Out_thrown_rData_branchInfo_0_predictPC;
  reg                 stage1Out_thrown_rData_branchInfo_0_predictResult;
  reg        [31:0]   stage1Out_thrown_rData_branchInfo_1_predictPC;
  reg                 stage1Out_thrown_rData_branchInfo_1_predictResult;
  reg                 stage1Out_thrown_rData_exceptionInfo_0_exception;
  reg        [5:0]    stage1Out_thrown_rData_exceptionInfo_0_eCode;
  reg        [0:0]    stage1Out_thrown_rData_exceptionInfo_0_eSubCode;
  reg                 stage1Out_thrown_rData_exceptionInfo_1_exception;
  reg        [5:0]    stage1Out_thrown_rData_exceptionInfo_1_eCode;
  reg        [0:0]    stage1Out_thrown_rData_exceptionInfo_1_eSubCode;
  reg        [31:0]   stage1Out_thrown_rData_pc_0;
  reg        [31:0]   stage1Out_thrown_rData_pc_1;
  reg        [1:0]    stage1Out_thrown_rData_valid;
  reg                 stage1Out_thrown_rData_tlb_hit;
  reg        [19:0]   stage1Out_thrown_rData_tlb_pageInfo_ppn;
  reg        [1:0]    stage1Out_thrown_rData_tlb_pageInfo_plv;
  reg        [1:0]    stage1Out_thrown_rData_tlb_pageInfo_mat;
  reg                 stage1Out_thrown_rData_tlb_pageInfo_d;
  reg                 stage1Out_thrown_rData_tlb_pageInfo_v;
  reg        [3:0]    stage1Out_thrown_rData_wayValid_0;
  reg        [3:0]    stage1Out_thrown_rData_wayValid_1;
  reg                 stage1Out_thrown_rData_isStoreTag;
  reg                 stage1Out_thrown_rData_isIndexInvalidate;
  reg                 stage1Out_thrown_rData_isHitInvalidate;
  wire                when_Stream_l369;
  reg        [1:0]    acceptMask;
  reg                 fetchMask_0;
  reg                 fetchMask_1;
  wire                stage1Out_fire;
  wire                _zz_io_output_availMask;
  wire                _zz_io_output_availMask_1;
  reg                 exceptionInfo1_0_exception;
  reg        [5:0]    exceptionInfo1_0_eCode;
  reg        [0:0]    exceptionInfo1_0_eSubCode;
  reg                 exceptionInfo1_1_exception;
  reg        [5:0]    exceptionInfo1_1_eCode;
  reg        [0:0]    exceptionInfo1_1_eSubCode;
  reg                 exceptionInfo2_exception;
  reg        [5:0]    exceptionInfo2_eCode;
  reg        [0:0]    exceptionInfo2_eSubCode;
  reg        [1:0]    availMask;
  wire       [1:0]    fireMask;
  reg        [1:0]    portAvail;
  wire       [31:0]   portData_0_inst;
  wire       [31:0]   portData_0_branchInfo_predictPC;
  wire                portData_0_branchInfo_predictResult;
  wire                portData_0_exceptionInfo_exception;
  wire       [5:0]    portData_0_exceptionInfo_eCode;
  wire       [0:0]    portData_0_exceptionInfo_eSubCode;
  wire       [31:0]   portData_0_pc;
  wire       [31:0]   portData_1_inst;
  wire       [31:0]   portData_1_branchInfo_predictPC;
  wire                portData_1_branchInfo_predictResult;
  wire                portData_1_exceptionInfo_exception;
  wire       [5:0]    portData_1_exceptionInfo_eCode;
  wire       [0:0]    portData_1_exceptionInfo_eSubCode;
  wire       [31:0]   portData_1_pc;
  reg        [1:0]    hasException;
  wire                when_Cache_l79;
  wire                when_Cache_l83;
  reg        [31:0]   missBuffer_0;
  reg        [31:0]   missBuffer_1;
  wire                _zz_missAddr;
  wire       [31:0]   missAddr;
  reg        [3:0]    replacingWay;
  reg        [5:0]    transferBlockOffset;
  reg        [5:0]    transferIndexOffset;
  reg        [19:0]   transferTag;
  reg                 transferUncached;
  wire       [31:0]   transferAddr;
  reg        [1:0]    sameBlockMask;
  reg        [1:0]    bufWriteMask;
  reg                 refilling;
  reg                 lruBit_0_0;
  reg                 lruBit_0_1;
  reg                 lruBit_0_2;
  reg                 lruBit_1_0;
  reg                 lruBit_1_1;
  reg                 lruBit_1_2;
  reg                 lruBit_2_0;
  reg                 lruBit_2_1;
  reg                 lruBit_2_2;
  reg                 lruBit_3_0;
  reg                 lruBit_3_1;
  reg                 lruBit_3_2;
  reg                 lruBit_4_0;
  reg                 lruBit_4_1;
  reg                 lruBit_4_2;
  reg                 lruBit_5_0;
  reg                 lruBit_5_1;
  reg                 lruBit_5_2;
  reg                 lruBit_6_0;
  reg                 lruBit_6_1;
  reg                 lruBit_6_2;
  reg                 lruBit_7_0;
  reg                 lruBit_7_1;
  reg                 lruBit_7_2;
  reg                 lruBit_8_0;
  reg                 lruBit_8_1;
  reg                 lruBit_8_2;
  reg                 lruBit_9_0;
  reg                 lruBit_9_1;
  reg                 lruBit_9_2;
  reg                 lruBit_10_0;
  reg                 lruBit_10_1;
  reg                 lruBit_10_2;
  reg                 lruBit_11_0;
  reg                 lruBit_11_1;
  reg                 lruBit_11_2;
  reg                 lruBit_12_0;
  reg                 lruBit_12_1;
  reg                 lruBit_12_2;
  reg                 lruBit_13_0;
  reg                 lruBit_13_1;
  reg                 lruBit_13_2;
  reg                 lruBit_14_0;
  reg                 lruBit_14_1;
  reg                 lruBit_14_2;
  reg                 lruBit_15_0;
  reg                 lruBit_15_1;
  reg                 lruBit_15_2;
  reg                 lruBit_16_0;
  reg                 lruBit_16_1;
  reg                 lruBit_16_2;
  reg                 lruBit_17_0;
  reg                 lruBit_17_1;
  reg                 lruBit_17_2;
  reg                 lruBit_18_0;
  reg                 lruBit_18_1;
  reg                 lruBit_18_2;
  reg                 lruBit_19_0;
  reg                 lruBit_19_1;
  reg                 lruBit_19_2;
  reg                 lruBit_20_0;
  reg                 lruBit_20_1;
  reg                 lruBit_20_2;
  reg                 lruBit_21_0;
  reg                 lruBit_21_1;
  reg                 lruBit_21_2;
  reg                 lruBit_22_0;
  reg                 lruBit_22_1;
  reg                 lruBit_22_2;
  reg                 lruBit_23_0;
  reg                 lruBit_23_1;
  reg                 lruBit_23_2;
  reg                 lruBit_24_0;
  reg                 lruBit_24_1;
  reg                 lruBit_24_2;
  reg                 lruBit_25_0;
  reg                 lruBit_25_1;
  reg                 lruBit_25_2;
  reg                 lruBit_26_0;
  reg                 lruBit_26_1;
  reg                 lruBit_26_2;
  reg                 lruBit_27_0;
  reg                 lruBit_27_1;
  reg                 lruBit_27_2;
  reg                 lruBit_28_0;
  reg                 lruBit_28_1;
  reg                 lruBit_28_2;
  reg                 lruBit_29_0;
  reg                 lruBit_29_1;
  reg                 lruBit_29_2;
  reg                 lruBit_30_0;
  reg                 lruBit_30_1;
  reg                 lruBit_30_2;
  reg                 lruBit_31_0;
  reg                 lruBit_31_1;
  reg                 lruBit_31_2;
  reg        [3:0]    wayToReplace_0;
  reg        [3:0]    wayToReplace_1;
  reg        [3:0]    wayOfReplace_0;
  reg        [3:0]    wayOfReplace_1;
  wire                when_Cache_l131;
  wire                when_Cache_l311;
  wire       [31:0]   _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                _zz_14;
  wire                _zz_15;
  wire                _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_lruBit_0_0;
  wire                when_Cache_l311_1;
  wire                _zz_lruBit_0_1;
  wire                when_Cache_l311_2;
  wire                _zz_lruBit_0_2;
  wire                when_Cache_l131_1;
  wire                when_Cache_l311_3;
  wire       [31:0]   _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire                _zz_lruBit_0_0_1;
  wire                when_Cache_l311_4;
  wire                _zz_lruBit_0_1_1;
  wire                when_Cache_l311_5;
  wire                _zz_lruBit_0_2_1;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg        [1:0]    allowMask;
  wire                when_Cache_l222;
  wire                io_input_0_fire;
  wire                _zz_portData_0_inst;
  wire                _zz_portData_0_inst_1;
  wire                _zz_portData_0_inst_2;
  wire                when_Cache_l255;
  wire       [0:0]    _zz_io_output_info_0_inst;
  reg        [1:0]    _zz_wayToReplace_0;
  reg        [1:0]    _zz_wayToReplace_0_1;
  reg        [1:0]    _zz_wayToReplace_0_2;
  reg        [1:0]    _zz_wayToReplace_0_3;
  wire                when_Cache_l222_1;
  wire                io_input_1_fire;
  wire                _zz_portData_1_inst;
  wire                _zz_portData_1_inst_1;
  wire                _zz_portData_1_inst_2;
  wire                when_Cache_l255_1;
  wire       [0:0]    _zz_io_output_info_1_inst;
  reg        [1:0]    _zz_wayToReplace_1;
  reg        [1:0]    _zz_wayToReplace_1_1;
  reg        [1:0]    _zz_wayToReplace_1_2;
  reg        [1:0]    _zz_wayToReplace_1_3;
  wire       [4:0]    cacopIdx;
  wire       [3:0]    cacopWay;
  wire                when_Cache_l283;
  wire                when_Cache_l285;
  wire       [31:0]   _zz_67;
  wire                when_Cache_l285_1;
  wire       [31:0]   _zz_68;
  wire                when_Cache_l285_2;
  wire       [31:0]   _zz_69;
  wire                when_Cache_l285_3;
  wire       [31:0]   _zz_70;
  reg        [1:0]    fsm_stateReg;
  reg        [1:0]    fsm_stateNext;
  wire                when_Cache_l158;
  wire                when_Cache_l174;
  wire                when_Cache_l198;
  wire                when_Cache_l200;
  wire                when_Cache_l201;
  wire       [8:0]    _zz_wr_addr;
  wire       [31:0]   _zz_wr_data;
  wire                when_Cache_l200_1;
  wire                when_Cache_l201_1;
  wire       [8:0]    _zz_wr_addr_1;
  wire       [31:0]   _zz_wr_data_1;
  wire                when_Cache_l200_2;
  wire                when_Cache_l201_2;
  wire       [8:0]    _zz_wr_addr_2;
  wire       [31:0]   _zz_wr_data_2;
  wire                when_Cache_l200_3;
  wire                when_Cache_l201_3;
  wire       [8:0]    _zz_wr_addr_3;
  wire       [31:0]   _zz_wr_data_3;
  wire                when_Cache_l209;
  wire                when_Cache_l210;
  wire                when_StateMachine_l253;
  wire                when_StateMachine_l253_1;
  wire                when_Cache_l180;
  wire                when_Cache_l182;
  wire       [4:0]    _zz_wr_addr_4;
  wire       [20:0]   _zz_wr_data_4;
  wire       [31:0]   _zz_71;
  wire                when_Cache_l182_1;
  wire       [4:0]    _zz_wr_addr_5;
  wire       [20:0]   _zz_wr_data_5;
  wire       [31:0]   _zz_72;
  wire                when_Cache_l182_2;
  wire       [4:0]    _zz_wr_addr_6;
  wire       [20:0]   _zz_wr_data_6;
  wire       [31:0]   _zz_73;
  wire                when_Cache_l182_3;
  wire       [4:0]    _zz_wr_addr_7;
  wire       [20:0]   _zz_wr_data_7;
  wire       [31:0]   _zz_74;
  wire                when_Cache_l188;
  wire                when_Cache_l188_1;
  `ifndef SYNTHESIS
  reg [63:0] io_input_0_payload_size_string;
  reg [63:0] io_input_1_payload_size_string;
  reg [31:0] fsm_stateReg_string;
  reg [31:0] fsm_stateNext_string;
  `endif


  assign _zz_acceptMask = (io_output_allowMask <<< _zz_acceptMask_1);
  assign _zz_stage1Out_payload_wayValid_0_2 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_hit_0_1 = 1'b1;
  assign _zz_hit_0 = {1'd0, _zz_hit_0_1};
  assign _zz_stage1Out_payload_wayValid_0_5 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_hit_0_3 = 1'b1;
  assign _zz_hit_0_2 = {1'd0, _zz_hit_0_3};
  assign _zz_stage1Out_payload_wayValid_0_8 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_hit_0_5 = 1'b1;
  assign _zz_hit_0_4 = {1'd0, _zz_hit_0_5};
  assign _zz_stage1Out_payload_wayValid_0_11 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_hit_0_7 = 1'b1;
  assign _zz_hit_0_6 = {1'd0, _zz_hit_0_7};
  assign _zz_hit_1_1 = 1'b1;
  assign _zz_hit_1 = {1'd0, _zz_hit_1_1};
  assign _zz_hit_1_3 = 1'b1;
  assign _zz_hit_1_2 = {1'd0, _zz_hit_1_3};
  assign _zz_hit_1_5 = 1'b1;
  assign _zz_hit_1_4 = {1'd0, _zz_hit_1_5};
  assign _zz_hit_1_7 = 1'b1;
  assign _zz_hit_1_6 = {1'd0, _zz_hit_1_7};
  assign _zz_exceptionInfo2_eCode = 2'b11;
  assign _zz_exceptionInfo2_eCode_1 = 3'b111;
  assign _zz_exceptionInfo2_eCode_2 = 3'b111;
  assign _zz_when_Cache_l131_1 = 1'b1;
  assign _zz_when_Cache_l131 = {1'd0, _zz_when_Cache_l131_1};
  assign _zz_when_Cache_l131_1_2 = 1'b1;
  assign _zz_when_Cache_l131_1_1 = {1'd0, _zz_when_Cache_l131_1_2};
  assign _zz_io_axi_arlen_1 = 4'b1111;
  assign _zz_io_axi_arlen = {4'd0, _zz_io_axi_arlen_1};
  assign _zz_exceptionInfo1_0_eCode = 4'b1000;
  assign _zz_exceptionInfo1_0_eCode_1 = 4'b1000;
  assign _zz__zz_io_output_info_0_inst = (2'b00 + _zz__zz_io_output_info_0_inst_1);
  assign _zz_exceptionInfo1_1_eCode = 4'b1000;
  assign _zz_exceptionInfo1_1_eCode_1 = 4'b1000;
  assign _zz__zz_io_output_info_1_inst = (2'b01 + _zz__zz_io_output_info_1_inst_1);
  assign _zz_cacopWay = (4'b0001 <<< stage2In_payload_pc_0[1 : 0]);
  assign _zz_when_Cache_l198_1 = 1'b1;
  assign _zz_when_Cache_l198 = {1'd0, _zz_when_Cache_l198_1};
  assign _zz_when_Cache_l180_1 = 1'b1;
  assign _zz_when_Cache_l180 = {1'd0, _zz_when_Cache_l180_1};
  assign _zz_rd_addr = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_rd_addr_1 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_rd_addr_2 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_rd_addr_3 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_rd_addr_4 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_rd_addr_5 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_rd_addr_6 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_rd_addr_7 = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign _zz_acceptMask_2 = {_zz_io_output_availMask_1,_zz_io_output_availMask};
  assign _zz_stage1Out_payload_wayValid_0_1 = _zz_stage1Out_payload_wayValid_0_2[10 : 6];
  assign _zz_stage1Out_payload_wayValid_0_4 = _zz_stage1Out_payload_wayValid_0_5[10 : 6];
  assign _zz_stage1Out_payload_wayValid_0_7 = _zz_stage1Out_payload_wayValid_0_8[10 : 6];
  assign _zz_stage1Out_payload_wayValid_0_10 = _zz_stage1Out_payload_wayValid_0_11[10 : 6];
  assign _zz_stage1Out_payload_wayValid_1_1 = io_input_1_payload_address[10 : 6];
  assign _zz_stage1Out_payload_wayValid_1_3 = io_input_1_payload_address[10 : 6];
  assign _zz_stage1Out_payload_wayValid_1_5 = io_input_1_payload_address[10 : 6];
  assign _zz_stage1Out_payload_wayValid_1_7 = io_input_1_payload_address[10 : 6];
  assign _zz_fireMask_1 = {_zz_io_output_availMask_1,_zz_io_output_availMask};
  assign _zz_portData_0_inst_4 = {_zz_portData_0_inst_2,_zz_portData_0_inst_1};
  assign _zz__zz_io_output_info_0_inst_2 = {_zz_io_output_availMask_1,_zz_io_output_availMask};
  assign _zz__zz_wayToReplace_0_1 = stage2In_payload_pc_0[10 : 6];
  assign _zz__zz_wayToReplace_0_3 = stage2In_payload_pc_0[10 : 6];
  assign _zz__zz_wayToReplace_0_1_2 = stage2In_payload_pc_0[10 : 6];
  assign _zz__zz_wayToReplace_0_1_4 = stage2In_payload_pc_0[10 : 6];
  assign _zz__zz_wayToReplace_0_2_2 = stage2In_payload_pc_0[10 : 6];
  assign _zz__zz_wayToReplace_0_2_4 = stage2In_payload_pc_0[10 : 6];
  assign _zz__zz_wayToReplace_0_3_2 = stage2In_payload_pc_0[10 : 6];
  assign _zz__zz_wayToReplace_0_3_4 = stage2In_payload_pc_0[10 : 6];
  assign _zz_portData_1_inst_4 = {_zz_portData_1_inst_2,_zz_portData_1_inst_1};
  assign _zz__zz_io_output_info_1_inst_2 = {_zz_io_output_availMask_1,_zz_io_output_availMask};
  assign _zz__zz_wayToReplace_1_1 = stage2In_payload_pc_1[10 : 6];
  assign _zz__zz_wayToReplace_1_3 = stage2In_payload_pc_1[10 : 6];
  assign _zz__zz_wayToReplace_1_1_2 = stage2In_payload_pc_1[10 : 6];
  assign _zz__zz_wayToReplace_1_1_4 = stage2In_payload_pc_1[10 : 6];
  assign _zz__zz_wayToReplace_1_2_2 = stage2In_payload_pc_1[10 : 6];
  assign _zz__zz_wayToReplace_1_2_4 = stage2In_payload_pc_1[10 : 6];
  assign _zz__zz_wayToReplace_1_3_2 = stage2In_payload_pc_1[10 : 6];
  assign _zz__zz_wayToReplace_1_3_4 = stage2In_payload_pc_1[10 : 6];
  assign _zz_io_output_availMask_3 = {_zz_io_output_availMask_1,_zz_io_output_availMask};
  Ram_1w_1rs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(9),
    .wrDataWidth(32),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(9),
    .rdDataWidth(32)
  ) data_0 (
    .wr_clk  (aclk                ), //i
    .wr_en   (data_0_wr_en        ), //i
    .wr_mask (data_0_wr_mask      ), //i
    .wr_addr (_zz_wr_addr[8:0]    ), //i
    .wr_data (_zz_wr_data[31:0]   ), //i
    .rd_clk  (aclk                ), //i
    .rd_en   (data_0_rd_en        ), //i
    .rd_addr (data_0_rd_addr[8:0] ), //i
    .rd_data (data_0_rd_data[31:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(9),
    .wrDataWidth(32),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(9),
    .rdDataWidth(32)
  ) data_0_1 (
    .wr_clk  (aclk                  ), //i
    .wr_en   (data_0_1_wr_en        ), //i
    .wr_mask (data_0_1_wr_mask      ), //i
    .wr_addr (_zz_wr_addr[8:0]      ), //i
    .wr_data (_zz_wr_data[31:0]     ), //i
    .rd_clk  (aclk                  ), //i
    .rd_en   (data_0_1_rd_en        ), //i
    .rd_addr (data_0_1_rd_addr[8:0] ), //i
    .rd_data (data_0_1_rd_data[31:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(9),
    .wrDataWidth(32),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(9),
    .rdDataWidth(32)
  ) data_1 (
    .wr_clk  (aclk                ), //i
    .wr_en   (data_1_wr_en        ), //i
    .wr_mask (data_1_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_1[8:0]  ), //i
    .wr_data (_zz_wr_data_1[31:0] ), //i
    .rd_clk  (aclk                ), //i
    .rd_en   (data_1_rd_en        ), //i
    .rd_addr (data_1_rd_addr[8:0] ), //i
    .rd_data (data_1_rd_data[31:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(9),
    .wrDataWidth(32),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(9),
    .rdDataWidth(32)
  ) data_1_1 (
    .wr_clk  (aclk                  ), //i
    .wr_en   (data_1_1_wr_en        ), //i
    .wr_mask (data_1_1_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_1[8:0]    ), //i
    .wr_data (_zz_wr_data_1[31:0]   ), //i
    .rd_clk  (aclk                  ), //i
    .rd_en   (data_1_1_rd_en        ), //i
    .rd_addr (data_1_1_rd_addr[8:0] ), //i
    .rd_data (data_1_1_rd_data[31:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(9),
    .wrDataWidth(32),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(9),
    .rdDataWidth(32)
  ) data_2 (
    .wr_clk  (aclk                ), //i
    .wr_en   (data_2_wr_en        ), //i
    .wr_mask (data_2_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_2[8:0]  ), //i
    .wr_data (_zz_wr_data_2[31:0] ), //i
    .rd_clk  (aclk                ), //i
    .rd_en   (data_2_rd_en        ), //i
    .rd_addr (data_2_rd_addr[8:0] ), //i
    .rd_data (data_2_rd_data[31:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(9),
    .wrDataWidth(32),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(9),
    .rdDataWidth(32)
  ) data_2_1 (
    .wr_clk  (aclk                  ), //i
    .wr_en   (data_2_1_wr_en        ), //i
    .wr_mask (data_2_1_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_2[8:0]    ), //i
    .wr_data (_zz_wr_data_2[31:0]   ), //i
    .rd_clk  (aclk                  ), //i
    .rd_en   (data_2_1_rd_en        ), //i
    .rd_addr (data_2_1_rd_addr[8:0] ), //i
    .rd_data (data_2_1_rd_data[31:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(9),
    .wrDataWidth(32),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(9),
    .rdDataWidth(32)
  ) data_3 (
    .wr_clk  (aclk                ), //i
    .wr_en   (data_3_wr_en        ), //i
    .wr_mask (data_3_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_3[8:0]  ), //i
    .wr_data (_zz_wr_data_3[31:0] ), //i
    .rd_clk  (aclk                ), //i
    .rd_en   (data_3_rd_en        ), //i
    .rd_addr (data_3_rd_addr[8:0] ), //i
    .rd_data (data_3_rd_data[31:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(512),
    .wordWidth(32),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(9),
    .wrDataWidth(32),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(9),
    .rdDataWidth(32)
  ) data_3_1 (
    .wr_clk  (aclk                  ), //i
    .wr_en   (data_3_1_wr_en        ), //i
    .wr_mask (data_3_1_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_3[8:0]    ), //i
    .wr_data (_zz_wr_data_3[31:0]   ), //i
    .rd_clk  (aclk                  ), //i
    .rd_en   (data_3_1_rd_en        ), //i
    .rd_addr (data_3_1_rd_addr[8:0] ), //i
    .rd_data (data_3_1_rd_data[31:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_0 (
    .wr_clk  (aclk               ), //i
    .wr_en   (tag_0_wr_en        ), //i
    .wr_mask (tag_0_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_4[4:0] ), //i
    .wr_data (_zz_wr_data_4[20:0]), //i
    .rd_clk  (aclk               ), //i
    .rd_en   (tag_0_rd_en        ), //i
    .rd_addr (tag_0_rd_addr[4:0] ), //i
    .rd_data (tag_0_rd_data[20:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_0_1 (
    .wr_clk  (aclk                 ), //i
    .wr_en   (tag_0_1_wr_en        ), //i
    .wr_mask (tag_0_1_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_4[4:0]   ), //i
    .wr_data (_zz_wr_data_4[20:0]  ), //i
    .rd_clk  (aclk                 ), //i
    .rd_en   (tag_0_1_rd_en        ), //i
    .rd_addr (tag_0_1_rd_addr[4:0] ), //i
    .rd_data (tag_0_1_rd_data[20:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_1 (
    .wr_clk  (aclk               ), //i
    .wr_en   (tag_1_wr_en        ), //i
    .wr_mask (tag_1_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_5[4:0] ), //i
    .wr_data (_zz_wr_data_5[20:0]), //i
    .rd_clk  (aclk               ), //i
    .rd_en   (tag_1_rd_en        ), //i
    .rd_addr (tag_1_rd_addr[4:0] ), //i
    .rd_data (tag_1_rd_data[20:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_1_1 (
    .wr_clk  (aclk                 ), //i
    .wr_en   (tag_1_1_wr_en        ), //i
    .wr_mask (tag_1_1_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_5[4:0]   ), //i
    .wr_data (_zz_wr_data_5[20:0]  ), //i
    .rd_clk  (aclk                 ), //i
    .rd_en   (tag_1_1_rd_en        ), //i
    .rd_addr (tag_1_1_rd_addr[4:0] ), //i
    .rd_data (tag_1_1_rd_data[20:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_2 (
    .wr_clk  (aclk               ), //i
    .wr_en   (tag_2_wr_en        ), //i
    .wr_mask (tag_2_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_6[4:0] ), //i
    .wr_data (_zz_wr_data_6[20:0]), //i
    .rd_clk  (aclk               ), //i
    .rd_en   (tag_2_rd_en        ), //i
    .rd_addr (tag_2_rd_addr[4:0] ), //i
    .rd_data (tag_2_rd_data[20:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_2_1 (
    .wr_clk  (aclk                 ), //i
    .wr_en   (tag_2_1_wr_en        ), //i
    .wr_mask (tag_2_1_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_6[4:0]   ), //i
    .wr_data (_zz_wr_data_6[20:0]  ), //i
    .rd_clk  (aclk                 ), //i
    .rd_en   (tag_2_1_rd_en        ), //i
    .rd_addr (tag_2_1_rd_addr[4:0] ), //i
    .rd_data (tag_2_1_rd_data[20:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_3 (
    .wr_clk  (aclk               ), //i
    .wr_en   (tag_3_wr_en        ), //i
    .wr_mask (tag_3_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_7[4:0] ), //i
    .wr_data (_zz_wr_data_7[20:0]), //i
    .rd_clk  (aclk               ), //i
    .rd_en   (tag_3_rd_en        ), //i
    .rd_addr (tag_3_rd_addr[4:0] ), //i
    .rd_data (tag_3_rd_data[20:0])  //o
  );
  Ram_1w_1rs #(
    .wordCount(32),
    .wordWidth(21),
    .clockCrossing(1'b0),
    .technology("auto"),
    .readUnderWrite("dontCare"),
    .wrAddressWidth(5),
    .wrDataWidth(21),
    .wrMaskWidth(1),
    .wrMaskEnable(1'b0),
    .rdAddressWidth(5),
    .rdDataWidth(21)
  ) tag_3_1 (
    .wr_clk  (aclk                 ), //i
    .wr_en   (tag_3_1_wr_en        ), //i
    .wr_mask (tag_3_1_wr_mask      ), //i
    .wr_addr (_zz_wr_addr_7[4:0]   ), //i
    .wr_data (_zz_wr_data_7[20:0]  ), //i
    .rd_clk  (aclk                 ), //i
    .rd_en   (tag_3_1_rd_en        ), //i
    .rd_addr (tag_3_1_rd_addr[4:0] ), //i
    .rd_data (tag_3_1_rd_data[20:0])  //o
  );
  always @(*) begin
    case(_zz_acceptMask_2)
      2'b00 : _zz_acceptMask_1 = 2'b00;
      2'b01 : _zz_acceptMask_1 = 2'b01;
      2'b10 : _zz_acceptMask_1 = 2'b01;
      default : _zz_acceptMask_1 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_0_1)
      5'b00000 : _zz_stage1Out_payload_wayValid_0 = valid_0_0;
      5'b00001 : _zz_stage1Out_payload_wayValid_0 = valid_0_1;
      5'b00010 : _zz_stage1Out_payload_wayValid_0 = valid_0_2;
      5'b00011 : _zz_stage1Out_payload_wayValid_0 = valid_0_3;
      5'b00100 : _zz_stage1Out_payload_wayValid_0 = valid_0_4;
      5'b00101 : _zz_stage1Out_payload_wayValid_0 = valid_0_5;
      5'b00110 : _zz_stage1Out_payload_wayValid_0 = valid_0_6;
      5'b00111 : _zz_stage1Out_payload_wayValid_0 = valid_0_7;
      5'b01000 : _zz_stage1Out_payload_wayValid_0 = valid_0_8;
      5'b01001 : _zz_stage1Out_payload_wayValid_0 = valid_0_9;
      5'b01010 : _zz_stage1Out_payload_wayValid_0 = valid_0_10;
      5'b01011 : _zz_stage1Out_payload_wayValid_0 = valid_0_11;
      5'b01100 : _zz_stage1Out_payload_wayValid_0 = valid_0_12;
      5'b01101 : _zz_stage1Out_payload_wayValid_0 = valid_0_13;
      5'b01110 : _zz_stage1Out_payload_wayValid_0 = valid_0_14;
      5'b01111 : _zz_stage1Out_payload_wayValid_0 = valid_0_15;
      5'b10000 : _zz_stage1Out_payload_wayValid_0 = valid_0_16;
      5'b10001 : _zz_stage1Out_payload_wayValid_0 = valid_0_17;
      5'b10010 : _zz_stage1Out_payload_wayValid_0 = valid_0_18;
      5'b10011 : _zz_stage1Out_payload_wayValid_0 = valid_0_19;
      5'b10100 : _zz_stage1Out_payload_wayValid_0 = valid_0_20;
      5'b10101 : _zz_stage1Out_payload_wayValid_0 = valid_0_21;
      5'b10110 : _zz_stage1Out_payload_wayValid_0 = valid_0_22;
      5'b10111 : _zz_stage1Out_payload_wayValid_0 = valid_0_23;
      5'b11000 : _zz_stage1Out_payload_wayValid_0 = valid_0_24;
      5'b11001 : _zz_stage1Out_payload_wayValid_0 = valid_0_25;
      5'b11010 : _zz_stage1Out_payload_wayValid_0 = valid_0_26;
      5'b11011 : _zz_stage1Out_payload_wayValid_0 = valid_0_27;
      5'b11100 : _zz_stage1Out_payload_wayValid_0 = valid_0_28;
      5'b11101 : _zz_stage1Out_payload_wayValid_0 = valid_0_29;
      5'b11110 : _zz_stage1Out_payload_wayValid_0 = valid_0_30;
      default : _zz_stage1Out_payload_wayValid_0 = valid_0_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_0_4)
      5'b00000 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_0;
      5'b00001 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_1;
      5'b00010 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_2;
      5'b00011 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_3;
      5'b00100 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_4;
      5'b00101 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_5;
      5'b00110 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_6;
      5'b00111 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_7;
      5'b01000 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_8;
      5'b01001 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_9;
      5'b01010 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_10;
      5'b01011 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_11;
      5'b01100 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_12;
      5'b01101 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_13;
      5'b01110 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_14;
      5'b01111 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_15;
      5'b10000 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_16;
      5'b10001 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_17;
      5'b10010 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_18;
      5'b10011 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_19;
      5'b10100 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_20;
      5'b10101 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_21;
      5'b10110 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_22;
      5'b10111 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_23;
      5'b11000 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_24;
      5'b11001 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_25;
      5'b11010 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_26;
      5'b11011 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_27;
      5'b11100 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_28;
      5'b11101 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_29;
      5'b11110 : _zz_stage1Out_payload_wayValid_0_3 = valid_1_30;
      default : _zz_stage1Out_payload_wayValid_0_3 = valid_1_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_0_7)
      5'b00000 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_0;
      5'b00001 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_1;
      5'b00010 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_2;
      5'b00011 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_3;
      5'b00100 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_4;
      5'b00101 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_5;
      5'b00110 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_6;
      5'b00111 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_7;
      5'b01000 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_8;
      5'b01001 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_9;
      5'b01010 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_10;
      5'b01011 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_11;
      5'b01100 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_12;
      5'b01101 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_13;
      5'b01110 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_14;
      5'b01111 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_15;
      5'b10000 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_16;
      5'b10001 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_17;
      5'b10010 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_18;
      5'b10011 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_19;
      5'b10100 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_20;
      5'b10101 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_21;
      5'b10110 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_22;
      5'b10111 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_23;
      5'b11000 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_24;
      5'b11001 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_25;
      5'b11010 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_26;
      5'b11011 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_27;
      5'b11100 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_28;
      5'b11101 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_29;
      5'b11110 : _zz_stage1Out_payload_wayValid_0_6 = valid_2_30;
      default : _zz_stage1Out_payload_wayValid_0_6 = valid_2_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_0_10)
      5'b00000 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_0;
      5'b00001 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_1;
      5'b00010 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_2;
      5'b00011 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_3;
      5'b00100 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_4;
      5'b00101 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_5;
      5'b00110 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_6;
      5'b00111 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_7;
      5'b01000 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_8;
      5'b01001 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_9;
      5'b01010 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_10;
      5'b01011 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_11;
      5'b01100 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_12;
      5'b01101 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_13;
      5'b01110 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_14;
      5'b01111 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_15;
      5'b10000 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_16;
      5'b10001 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_17;
      5'b10010 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_18;
      5'b10011 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_19;
      5'b10100 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_20;
      5'b10101 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_21;
      5'b10110 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_22;
      5'b10111 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_23;
      5'b11000 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_24;
      5'b11001 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_25;
      5'b11010 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_26;
      5'b11011 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_27;
      5'b11100 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_28;
      5'b11101 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_29;
      5'b11110 : _zz_stage1Out_payload_wayValid_0_9 = valid_3_30;
      default : _zz_stage1Out_payload_wayValid_0_9 = valid_3_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_1_1)
      5'b00000 : _zz_stage1Out_payload_wayValid_1 = valid_0_0;
      5'b00001 : _zz_stage1Out_payload_wayValid_1 = valid_0_1;
      5'b00010 : _zz_stage1Out_payload_wayValid_1 = valid_0_2;
      5'b00011 : _zz_stage1Out_payload_wayValid_1 = valid_0_3;
      5'b00100 : _zz_stage1Out_payload_wayValid_1 = valid_0_4;
      5'b00101 : _zz_stage1Out_payload_wayValid_1 = valid_0_5;
      5'b00110 : _zz_stage1Out_payload_wayValid_1 = valid_0_6;
      5'b00111 : _zz_stage1Out_payload_wayValid_1 = valid_0_7;
      5'b01000 : _zz_stage1Out_payload_wayValid_1 = valid_0_8;
      5'b01001 : _zz_stage1Out_payload_wayValid_1 = valid_0_9;
      5'b01010 : _zz_stage1Out_payload_wayValid_1 = valid_0_10;
      5'b01011 : _zz_stage1Out_payload_wayValid_1 = valid_0_11;
      5'b01100 : _zz_stage1Out_payload_wayValid_1 = valid_0_12;
      5'b01101 : _zz_stage1Out_payload_wayValid_1 = valid_0_13;
      5'b01110 : _zz_stage1Out_payload_wayValid_1 = valid_0_14;
      5'b01111 : _zz_stage1Out_payload_wayValid_1 = valid_0_15;
      5'b10000 : _zz_stage1Out_payload_wayValid_1 = valid_0_16;
      5'b10001 : _zz_stage1Out_payload_wayValid_1 = valid_0_17;
      5'b10010 : _zz_stage1Out_payload_wayValid_1 = valid_0_18;
      5'b10011 : _zz_stage1Out_payload_wayValid_1 = valid_0_19;
      5'b10100 : _zz_stage1Out_payload_wayValid_1 = valid_0_20;
      5'b10101 : _zz_stage1Out_payload_wayValid_1 = valid_0_21;
      5'b10110 : _zz_stage1Out_payload_wayValid_1 = valid_0_22;
      5'b10111 : _zz_stage1Out_payload_wayValid_1 = valid_0_23;
      5'b11000 : _zz_stage1Out_payload_wayValid_1 = valid_0_24;
      5'b11001 : _zz_stage1Out_payload_wayValid_1 = valid_0_25;
      5'b11010 : _zz_stage1Out_payload_wayValid_1 = valid_0_26;
      5'b11011 : _zz_stage1Out_payload_wayValid_1 = valid_0_27;
      5'b11100 : _zz_stage1Out_payload_wayValid_1 = valid_0_28;
      5'b11101 : _zz_stage1Out_payload_wayValid_1 = valid_0_29;
      5'b11110 : _zz_stage1Out_payload_wayValid_1 = valid_0_30;
      default : _zz_stage1Out_payload_wayValid_1 = valid_0_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_1_3)
      5'b00000 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_0;
      5'b00001 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_1;
      5'b00010 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_2;
      5'b00011 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_3;
      5'b00100 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_4;
      5'b00101 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_5;
      5'b00110 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_6;
      5'b00111 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_7;
      5'b01000 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_8;
      5'b01001 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_9;
      5'b01010 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_10;
      5'b01011 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_11;
      5'b01100 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_12;
      5'b01101 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_13;
      5'b01110 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_14;
      5'b01111 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_15;
      5'b10000 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_16;
      5'b10001 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_17;
      5'b10010 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_18;
      5'b10011 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_19;
      5'b10100 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_20;
      5'b10101 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_21;
      5'b10110 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_22;
      5'b10111 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_23;
      5'b11000 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_24;
      5'b11001 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_25;
      5'b11010 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_26;
      5'b11011 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_27;
      5'b11100 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_28;
      5'b11101 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_29;
      5'b11110 : _zz_stage1Out_payload_wayValid_1_2 = valid_1_30;
      default : _zz_stage1Out_payload_wayValid_1_2 = valid_1_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_1_5)
      5'b00000 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_0;
      5'b00001 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_1;
      5'b00010 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_2;
      5'b00011 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_3;
      5'b00100 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_4;
      5'b00101 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_5;
      5'b00110 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_6;
      5'b00111 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_7;
      5'b01000 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_8;
      5'b01001 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_9;
      5'b01010 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_10;
      5'b01011 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_11;
      5'b01100 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_12;
      5'b01101 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_13;
      5'b01110 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_14;
      5'b01111 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_15;
      5'b10000 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_16;
      5'b10001 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_17;
      5'b10010 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_18;
      5'b10011 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_19;
      5'b10100 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_20;
      5'b10101 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_21;
      5'b10110 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_22;
      5'b10111 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_23;
      5'b11000 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_24;
      5'b11001 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_25;
      5'b11010 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_26;
      5'b11011 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_27;
      5'b11100 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_28;
      5'b11101 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_29;
      5'b11110 : _zz_stage1Out_payload_wayValid_1_4 = valid_2_30;
      default : _zz_stage1Out_payload_wayValid_1_4 = valid_2_31;
    endcase
  end

  always @(*) begin
    case(_zz_stage1Out_payload_wayValid_1_7)
      5'b00000 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_0;
      5'b00001 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_1;
      5'b00010 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_2;
      5'b00011 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_3;
      5'b00100 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_4;
      5'b00101 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_5;
      5'b00110 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_6;
      5'b00111 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_7;
      5'b01000 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_8;
      5'b01001 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_9;
      5'b01010 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_10;
      5'b01011 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_11;
      5'b01100 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_12;
      5'b01101 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_13;
      5'b01110 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_14;
      5'b01111 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_15;
      5'b10000 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_16;
      5'b10001 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_17;
      5'b10010 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_18;
      5'b10011 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_19;
      5'b10100 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_20;
      5'b10101 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_21;
      5'b10110 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_22;
      5'b10111 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_23;
      5'b11000 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_24;
      5'b11001 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_25;
      5'b11010 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_26;
      5'b11011 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_27;
      5'b11100 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_28;
      5'b11101 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_29;
      5'b11110 : _zz_stage1Out_payload_wayValid_1_6 = valid_3_30;
      default : _zz_stage1Out_payload_wayValid_1_6 = valid_3_31;
    endcase
  end

  always @(*) begin
    case(_zz_fireMask_1)
      2'b00 : _zz_fireMask = 2'b00;
      2'b01 : _zz_fireMask = 2'b01;
      2'b10 : _zz_fireMask = 2'b01;
      default : _zz_fireMask = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_portData_0_inst_4)
      2'b00 : _zz_portData_0_inst_3 = dataRead_0_0;
      2'b01 : _zz_portData_0_inst_3 = dataRead_0_1;
      2'b10 : _zz_portData_0_inst_3 = dataRead_0_2;
      default : _zz_portData_0_inst_3 = dataRead_0_3;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_output_info_0_inst_2)
      2'b00 : _zz__zz_io_output_info_0_inst_1 = 2'b00;
      2'b01 : _zz__zz_io_output_info_0_inst_1 = 2'b01;
      2'b10 : _zz__zz_io_output_info_0_inst_1 = 2'b01;
      default : _zz__zz_io_output_info_0_inst_1 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_io_output_info_0_inst)
      1'b0 : begin
        _zz_io_output_info_0_inst_1 = portData_0_inst;
        _zz_io_output_info_0_branchInfo_predictPC = portData_0_branchInfo_predictPC;
        _zz_io_output_info_0_branchInfo_predictResult = portData_0_branchInfo_predictResult;
        _zz_io_output_info_0_exceptionInfo_exception = portData_0_exceptionInfo_exception;
        _zz_io_output_info_0_exceptionInfo_eCode = portData_0_exceptionInfo_eCode;
        _zz_io_output_info_0_exceptionInfo_eSubCode = portData_0_exceptionInfo_eSubCode;
        _zz_io_output_info_0_pc = portData_0_pc;
      end
      default : begin
        _zz_io_output_info_0_inst_1 = portData_1_inst;
        _zz_io_output_info_0_branchInfo_predictPC = portData_1_branchInfo_predictPC;
        _zz_io_output_info_0_branchInfo_predictResult = portData_1_branchInfo_predictResult;
        _zz_io_output_info_0_exceptionInfo_exception = portData_1_exceptionInfo_exception;
        _zz_io_output_info_0_exceptionInfo_eCode = portData_1_exceptionInfo_eCode;
        _zz_io_output_info_0_exceptionInfo_eSubCode = portData_1_exceptionInfo_eSubCode;
        _zz_io_output_info_0_pc = portData_1_pc;
      end
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_0_1)
      5'b00000 : _zz__zz_wayToReplace_0 = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace_0 = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace_0 = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace_0 = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace_0 = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace_0 = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace_0 = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace_0 = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace_0 = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace_0 = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace_0 = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace_0 = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace_0 = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace_0 = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace_0 = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace_0 = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace_0 = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace_0 = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace_0 = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace_0 = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace_0 = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace_0 = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace_0 = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace_0 = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace_0 = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace_0 = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace_0 = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace_0 = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace_0 = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace_0 = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace_0 = lruBit_30_0;
      default : _zz__zz_wayToReplace_0 = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_0_3)
      5'b00000 : _zz__zz_wayToReplace_0_2 = lruBit_0_1;
      5'b00001 : _zz__zz_wayToReplace_0_2 = lruBit_1_1;
      5'b00010 : _zz__zz_wayToReplace_0_2 = lruBit_2_1;
      5'b00011 : _zz__zz_wayToReplace_0_2 = lruBit_3_1;
      5'b00100 : _zz__zz_wayToReplace_0_2 = lruBit_4_1;
      5'b00101 : _zz__zz_wayToReplace_0_2 = lruBit_5_1;
      5'b00110 : _zz__zz_wayToReplace_0_2 = lruBit_6_1;
      5'b00111 : _zz__zz_wayToReplace_0_2 = lruBit_7_1;
      5'b01000 : _zz__zz_wayToReplace_0_2 = lruBit_8_1;
      5'b01001 : _zz__zz_wayToReplace_0_2 = lruBit_9_1;
      5'b01010 : _zz__zz_wayToReplace_0_2 = lruBit_10_1;
      5'b01011 : _zz__zz_wayToReplace_0_2 = lruBit_11_1;
      5'b01100 : _zz__zz_wayToReplace_0_2 = lruBit_12_1;
      5'b01101 : _zz__zz_wayToReplace_0_2 = lruBit_13_1;
      5'b01110 : _zz__zz_wayToReplace_0_2 = lruBit_14_1;
      5'b01111 : _zz__zz_wayToReplace_0_2 = lruBit_15_1;
      5'b10000 : _zz__zz_wayToReplace_0_2 = lruBit_16_1;
      5'b10001 : _zz__zz_wayToReplace_0_2 = lruBit_17_1;
      5'b10010 : _zz__zz_wayToReplace_0_2 = lruBit_18_1;
      5'b10011 : _zz__zz_wayToReplace_0_2 = lruBit_19_1;
      5'b10100 : _zz__zz_wayToReplace_0_2 = lruBit_20_1;
      5'b10101 : _zz__zz_wayToReplace_0_2 = lruBit_21_1;
      5'b10110 : _zz__zz_wayToReplace_0_2 = lruBit_22_1;
      5'b10111 : _zz__zz_wayToReplace_0_2 = lruBit_23_1;
      5'b11000 : _zz__zz_wayToReplace_0_2 = lruBit_24_1;
      5'b11001 : _zz__zz_wayToReplace_0_2 = lruBit_25_1;
      5'b11010 : _zz__zz_wayToReplace_0_2 = lruBit_26_1;
      5'b11011 : _zz__zz_wayToReplace_0_2 = lruBit_27_1;
      5'b11100 : _zz__zz_wayToReplace_0_2 = lruBit_28_1;
      5'b11101 : _zz__zz_wayToReplace_0_2 = lruBit_29_1;
      5'b11110 : _zz__zz_wayToReplace_0_2 = lruBit_30_1;
      default : _zz__zz_wayToReplace_0_2 = lruBit_31_1;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_0_1_2)
      5'b00000 : _zz__zz_wayToReplace_0_1_1 = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace_0_1_1 = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace_0_1_1 = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace_0_1_1 = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace_0_1_1 = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace_0_1_1 = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace_0_1_1 = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace_0_1_1 = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace_0_1_1 = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace_0_1_1 = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace_0_1_1 = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace_0_1_1 = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace_0_1_1 = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace_0_1_1 = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace_0_1_1 = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace_0_1_1 = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace_0_1_1 = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace_0_1_1 = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace_0_1_1 = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace_0_1_1 = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace_0_1_1 = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace_0_1_1 = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace_0_1_1 = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace_0_1_1 = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace_0_1_1 = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace_0_1_1 = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace_0_1_1 = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace_0_1_1 = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace_0_1_1 = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace_0_1_1 = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace_0_1_1 = lruBit_30_0;
      default : _zz__zz_wayToReplace_0_1_1 = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_0_1_4)
      5'b00000 : _zz__zz_wayToReplace_0_1_3 = lruBit_0_1;
      5'b00001 : _zz__zz_wayToReplace_0_1_3 = lruBit_1_1;
      5'b00010 : _zz__zz_wayToReplace_0_1_3 = lruBit_2_1;
      5'b00011 : _zz__zz_wayToReplace_0_1_3 = lruBit_3_1;
      5'b00100 : _zz__zz_wayToReplace_0_1_3 = lruBit_4_1;
      5'b00101 : _zz__zz_wayToReplace_0_1_3 = lruBit_5_1;
      5'b00110 : _zz__zz_wayToReplace_0_1_3 = lruBit_6_1;
      5'b00111 : _zz__zz_wayToReplace_0_1_3 = lruBit_7_1;
      5'b01000 : _zz__zz_wayToReplace_0_1_3 = lruBit_8_1;
      5'b01001 : _zz__zz_wayToReplace_0_1_3 = lruBit_9_1;
      5'b01010 : _zz__zz_wayToReplace_0_1_3 = lruBit_10_1;
      5'b01011 : _zz__zz_wayToReplace_0_1_3 = lruBit_11_1;
      5'b01100 : _zz__zz_wayToReplace_0_1_3 = lruBit_12_1;
      5'b01101 : _zz__zz_wayToReplace_0_1_3 = lruBit_13_1;
      5'b01110 : _zz__zz_wayToReplace_0_1_3 = lruBit_14_1;
      5'b01111 : _zz__zz_wayToReplace_0_1_3 = lruBit_15_1;
      5'b10000 : _zz__zz_wayToReplace_0_1_3 = lruBit_16_1;
      5'b10001 : _zz__zz_wayToReplace_0_1_3 = lruBit_17_1;
      5'b10010 : _zz__zz_wayToReplace_0_1_3 = lruBit_18_1;
      5'b10011 : _zz__zz_wayToReplace_0_1_3 = lruBit_19_1;
      5'b10100 : _zz__zz_wayToReplace_0_1_3 = lruBit_20_1;
      5'b10101 : _zz__zz_wayToReplace_0_1_3 = lruBit_21_1;
      5'b10110 : _zz__zz_wayToReplace_0_1_3 = lruBit_22_1;
      5'b10111 : _zz__zz_wayToReplace_0_1_3 = lruBit_23_1;
      5'b11000 : _zz__zz_wayToReplace_0_1_3 = lruBit_24_1;
      5'b11001 : _zz__zz_wayToReplace_0_1_3 = lruBit_25_1;
      5'b11010 : _zz__zz_wayToReplace_0_1_3 = lruBit_26_1;
      5'b11011 : _zz__zz_wayToReplace_0_1_3 = lruBit_27_1;
      5'b11100 : _zz__zz_wayToReplace_0_1_3 = lruBit_28_1;
      5'b11101 : _zz__zz_wayToReplace_0_1_3 = lruBit_29_1;
      5'b11110 : _zz__zz_wayToReplace_0_1_3 = lruBit_30_1;
      default : _zz__zz_wayToReplace_0_1_3 = lruBit_31_1;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_0_2_2)
      5'b00000 : _zz__zz_wayToReplace_0_2_1 = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace_0_2_1 = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace_0_2_1 = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace_0_2_1 = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace_0_2_1 = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace_0_2_1 = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace_0_2_1 = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace_0_2_1 = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace_0_2_1 = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace_0_2_1 = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace_0_2_1 = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace_0_2_1 = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace_0_2_1 = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace_0_2_1 = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace_0_2_1 = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace_0_2_1 = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace_0_2_1 = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace_0_2_1 = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace_0_2_1 = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace_0_2_1 = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace_0_2_1 = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace_0_2_1 = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace_0_2_1 = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace_0_2_1 = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace_0_2_1 = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace_0_2_1 = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace_0_2_1 = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace_0_2_1 = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace_0_2_1 = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace_0_2_1 = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace_0_2_1 = lruBit_30_0;
      default : _zz__zz_wayToReplace_0_2_1 = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_0_2_4)
      5'b00000 : _zz__zz_wayToReplace_0_2_3 = lruBit_0_2;
      5'b00001 : _zz__zz_wayToReplace_0_2_3 = lruBit_1_2;
      5'b00010 : _zz__zz_wayToReplace_0_2_3 = lruBit_2_2;
      5'b00011 : _zz__zz_wayToReplace_0_2_3 = lruBit_3_2;
      5'b00100 : _zz__zz_wayToReplace_0_2_3 = lruBit_4_2;
      5'b00101 : _zz__zz_wayToReplace_0_2_3 = lruBit_5_2;
      5'b00110 : _zz__zz_wayToReplace_0_2_3 = lruBit_6_2;
      5'b00111 : _zz__zz_wayToReplace_0_2_3 = lruBit_7_2;
      5'b01000 : _zz__zz_wayToReplace_0_2_3 = lruBit_8_2;
      5'b01001 : _zz__zz_wayToReplace_0_2_3 = lruBit_9_2;
      5'b01010 : _zz__zz_wayToReplace_0_2_3 = lruBit_10_2;
      5'b01011 : _zz__zz_wayToReplace_0_2_3 = lruBit_11_2;
      5'b01100 : _zz__zz_wayToReplace_0_2_3 = lruBit_12_2;
      5'b01101 : _zz__zz_wayToReplace_0_2_3 = lruBit_13_2;
      5'b01110 : _zz__zz_wayToReplace_0_2_3 = lruBit_14_2;
      5'b01111 : _zz__zz_wayToReplace_0_2_3 = lruBit_15_2;
      5'b10000 : _zz__zz_wayToReplace_0_2_3 = lruBit_16_2;
      5'b10001 : _zz__zz_wayToReplace_0_2_3 = lruBit_17_2;
      5'b10010 : _zz__zz_wayToReplace_0_2_3 = lruBit_18_2;
      5'b10011 : _zz__zz_wayToReplace_0_2_3 = lruBit_19_2;
      5'b10100 : _zz__zz_wayToReplace_0_2_3 = lruBit_20_2;
      5'b10101 : _zz__zz_wayToReplace_0_2_3 = lruBit_21_2;
      5'b10110 : _zz__zz_wayToReplace_0_2_3 = lruBit_22_2;
      5'b10111 : _zz__zz_wayToReplace_0_2_3 = lruBit_23_2;
      5'b11000 : _zz__zz_wayToReplace_0_2_3 = lruBit_24_2;
      5'b11001 : _zz__zz_wayToReplace_0_2_3 = lruBit_25_2;
      5'b11010 : _zz__zz_wayToReplace_0_2_3 = lruBit_26_2;
      5'b11011 : _zz__zz_wayToReplace_0_2_3 = lruBit_27_2;
      5'b11100 : _zz__zz_wayToReplace_0_2_3 = lruBit_28_2;
      5'b11101 : _zz__zz_wayToReplace_0_2_3 = lruBit_29_2;
      5'b11110 : _zz__zz_wayToReplace_0_2_3 = lruBit_30_2;
      default : _zz__zz_wayToReplace_0_2_3 = lruBit_31_2;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_0_3_2)
      5'b00000 : _zz__zz_wayToReplace_0_3_1 = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace_0_3_1 = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace_0_3_1 = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace_0_3_1 = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace_0_3_1 = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace_0_3_1 = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace_0_3_1 = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace_0_3_1 = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace_0_3_1 = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace_0_3_1 = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace_0_3_1 = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace_0_3_1 = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace_0_3_1 = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace_0_3_1 = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace_0_3_1 = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace_0_3_1 = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace_0_3_1 = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace_0_3_1 = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace_0_3_1 = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace_0_3_1 = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace_0_3_1 = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace_0_3_1 = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace_0_3_1 = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace_0_3_1 = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace_0_3_1 = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace_0_3_1 = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace_0_3_1 = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace_0_3_1 = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace_0_3_1 = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace_0_3_1 = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace_0_3_1 = lruBit_30_0;
      default : _zz__zz_wayToReplace_0_3_1 = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_0_3_4)
      5'b00000 : _zz__zz_wayToReplace_0_3_3 = lruBit_0_2;
      5'b00001 : _zz__zz_wayToReplace_0_3_3 = lruBit_1_2;
      5'b00010 : _zz__zz_wayToReplace_0_3_3 = lruBit_2_2;
      5'b00011 : _zz__zz_wayToReplace_0_3_3 = lruBit_3_2;
      5'b00100 : _zz__zz_wayToReplace_0_3_3 = lruBit_4_2;
      5'b00101 : _zz__zz_wayToReplace_0_3_3 = lruBit_5_2;
      5'b00110 : _zz__zz_wayToReplace_0_3_3 = lruBit_6_2;
      5'b00111 : _zz__zz_wayToReplace_0_3_3 = lruBit_7_2;
      5'b01000 : _zz__zz_wayToReplace_0_3_3 = lruBit_8_2;
      5'b01001 : _zz__zz_wayToReplace_0_3_3 = lruBit_9_2;
      5'b01010 : _zz__zz_wayToReplace_0_3_3 = lruBit_10_2;
      5'b01011 : _zz__zz_wayToReplace_0_3_3 = lruBit_11_2;
      5'b01100 : _zz__zz_wayToReplace_0_3_3 = lruBit_12_2;
      5'b01101 : _zz__zz_wayToReplace_0_3_3 = lruBit_13_2;
      5'b01110 : _zz__zz_wayToReplace_0_3_3 = lruBit_14_2;
      5'b01111 : _zz__zz_wayToReplace_0_3_3 = lruBit_15_2;
      5'b10000 : _zz__zz_wayToReplace_0_3_3 = lruBit_16_2;
      5'b10001 : _zz__zz_wayToReplace_0_3_3 = lruBit_17_2;
      5'b10010 : _zz__zz_wayToReplace_0_3_3 = lruBit_18_2;
      5'b10011 : _zz__zz_wayToReplace_0_3_3 = lruBit_19_2;
      5'b10100 : _zz__zz_wayToReplace_0_3_3 = lruBit_20_2;
      5'b10101 : _zz__zz_wayToReplace_0_3_3 = lruBit_21_2;
      5'b10110 : _zz__zz_wayToReplace_0_3_3 = lruBit_22_2;
      5'b10111 : _zz__zz_wayToReplace_0_3_3 = lruBit_23_2;
      5'b11000 : _zz__zz_wayToReplace_0_3_3 = lruBit_24_2;
      5'b11001 : _zz__zz_wayToReplace_0_3_3 = lruBit_25_2;
      5'b11010 : _zz__zz_wayToReplace_0_3_3 = lruBit_26_2;
      5'b11011 : _zz__zz_wayToReplace_0_3_3 = lruBit_27_2;
      5'b11100 : _zz__zz_wayToReplace_0_3_3 = lruBit_28_2;
      5'b11101 : _zz__zz_wayToReplace_0_3_3 = lruBit_29_2;
      5'b11110 : _zz__zz_wayToReplace_0_3_3 = lruBit_30_2;
      default : _zz__zz_wayToReplace_0_3_3 = lruBit_31_2;
    endcase
  end

  always @(*) begin
    case(_zz_portData_1_inst_4)
      2'b00 : _zz_portData_1_inst_3 = dataRead_1_0;
      2'b01 : _zz_portData_1_inst_3 = dataRead_1_1;
      2'b10 : _zz_portData_1_inst_3 = dataRead_1_2;
      default : _zz_portData_1_inst_3 = dataRead_1_3;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_output_info_1_inst_2)
      2'b00 : _zz__zz_io_output_info_1_inst_1 = 2'b00;
      2'b01 : _zz__zz_io_output_info_1_inst_1 = 2'b01;
      2'b10 : _zz__zz_io_output_info_1_inst_1 = 2'b01;
      default : _zz__zz_io_output_info_1_inst_1 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_io_output_info_1_inst)
      1'b0 : begin
        _zz_io_output_info_1_inst_1 = portData_0_inst;
        _zz_io_output_info_1_branchInfo_predictPC = portData_0_branchInfo_predictPC;
        _zz_io_output_info_1_branchInfo_predictResult = portData_0_branchInfo_predictResult;
        _zz_io_output_info_1_exceptionInfo_exception = portData_0_exceptionInfo_exception;
        _zz_io_output_info_1_exceptionInfo_eCode = portData_0_exceptionInfo_eCode;
        _zz_io_output_info_1_exceptionInfo_eSubCode = portData_0_exceptionInfo_eSubCode;
        _zz_io_output_info_1_pc = portData_0_pc;
      end
      default : begin
        _zz_io_output_info_1_inst_1 = portData_1_inst;
        _zz_io_output_info_1_branchInfo_predictPC = portData_1_branchInfo_predictPC;
        _zz_io_output_info_1_branchInfo_predictResult = portData_1_branchInfo_predictResult;
        _zz_io_output_info_1_exceptionInfo_exception = portData_1_exceptionInfo_exception;
        _zz_io_output_info_1_exceptionInfo_eCode = portData_1_exceptionInfo_eCode;
        _zz_io_output_info_1_exceptionInfo_eSubCode = portData_1_exceptionInfo_eSubCode;
        _zz_io_output_info_1_pc = portData_1_pc;
      end
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_1_1)
      5'b00000 : _zz__zz_wayToReplace_1 = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace_1 = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace_1 = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace_1 = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace_1 = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace_1 = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace_1 = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace_1 = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace_1 = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace_1 = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace_1 = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace_1 = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace_1 = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace_1 = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace_1 = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace_1 = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace_1 = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace_1 = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace_1 = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace_1 = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace_1 = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace_1 = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace_1 = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace_1 = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace_1 = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace_1 = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace_1 = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace_1 = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace_1 = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace_1 = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace_1 = lruBit_30_0;
      default : _zz__zz_wayToReplace_1 = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_1_3)
      5'b00000 : _zz__zz_wayToReplace_1_2 = lruBit_0_1;
      5'b00001 : _zz__zz_wayToReplace_1_2 = lruBit_1_1;
      5'b00010 : _zz__zz_wayToReplace_1_2 = lruBit_2_1;
      5'b00011 : _zz__zz_wayToReplace_1_2 = lruBit_3_1;
      5'b00100 : _zz__zz_wayToReplace_1_2 = lruBit_4_1;
      5'b00101 : _zz__zz_wayToReplace_1_2 = lruBit_5_1;
      5'b00110 : _zz__zz_wayToReplace_1_2 = lruBit_6_1;
      5'b00111 : _zz__zz_wayToReplace_1_2 = lruBit_7_1;
      5'b01000 : _zz__zz_wayToReplace_1_2 = lruBit_8_1;
      5'b01001 : _zz__zz_wayToReplace_1_2 = lruBit_9_1;
      5'b01010 : _zz__zz_wayToReplace_1_2 = lruBit_10_1;
      5'b01011 : _zz__zz_wayToReplace_1_2 = lruBit_11_1;
      5'b01100 : _zz__zz_wayToReplace_1_2 = lruBit_12_1;
      5'b01101 : _zz__zz_wayToReplace_1_2 = lruBit_13_1;
      5'b01110 : _zz__zz_wayToReplace_1_2 = lruBit_14_1;
      5'b01111 : _zz__zz_wayToReplace_1_2 = lruBit_15_1;
      5'b10000 : _zz__zz_wayToReplace_1_2 = lruBit_16_1;
      5'b10001 : _zz__zz_wayToReplace_1_2 = lruBit_17_1;
      5'b10010 : _zz__zz_wayToReplace_1_2 = lruBit_18_1;
      5'b10011 : _zz__zz_wayToReplace_1_2 = lruBit_19_1;
      5'b10100 : _zz__zz_wayToReplace_1_2 = lruBit_20_1;
      5'b10101 : _zz__zz_wayToReplace_1_2 = lruBit_21_1;
      5'b10110 : _zz__zz_wayToReplace_1_2 = lruBit_22_1;
      5'b10111 : _zz__zz_wayToReplace_1_2 = lruBit_23_1;
      5'b11000 : _zz__zz_wayToReplace_1_2 = lruBit_24_1;
      5'b11001 : _zz__zz_wayToReplace_1_2 = lruBit_25_1;
      5'b11010 : _zz__zz_wayToReplace_1_2 = lruBit_26_1;
      5'b11011 : _zz__zz_wayToReplace_1_2 = lruBit_27_1;
      5'b11100 : _zz__zz_wayToReplace_1_2 = lruBit_28_1;
      5'b11101 : _zz__zz_wayToReplace_1_2 = lruBit_29_1;
      5'b11110 : _zz__zz_wayToReplace_1_2 = lruBit_30_1;
      default : _zz__zz_wayToReplace_1_2 = lruBit_31_1;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_1_1_2)
      5'b00000 : _zz__zz_wayToReplace_1_1_1 = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace_1_1_1 = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace_1_1_1 = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace_1_1_1 = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace_1_1_1 = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace_1_1_1 = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace_1_1_1 = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace_1_1_1 = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace_1_1_1 = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace_1_1_1 = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace_1_1_1 = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace_1_1_1 = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace_1_1_1 = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace_1_1_1 = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace_1_1_1 = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace_1_1_1 = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace_1_1_1 = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace_1_1_1 = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace_1_1_1 = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace_1_1_1 = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace_1_1_1 = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace_1_1_1 = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace_1_1_1 = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace_1_1_1 = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace_1_1_1 = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace_1_1_1 = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace_1_1_1 = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace_1_1_1 = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace_1_1_1 = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace_1_1_1 = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace_1_1_1 = lruBit_30_0;
      default : _zz__zz_wayToReplace_1_1_1 = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_1_1_4)
      5'b00000 : _zz__zz_wayToReplace_1_1_3 = lruBit_0_1;
      5'b00001 : _zz__zz_wayToReplace_1_1_3 = lruBit_1_1;
      5'b00010 : _zz__zz_wayToReplace_1_1_3 = lruBit_2_1;
      5'b00011 : _zz__zz_wayToReplace_1_1_3 = lruBit_3_1;
      5'b00100 : _zz__zz_wayToReplace_1_1_3 = lruBit_4_1;
      5'b00101 : _zz__zz_wayToReplace_1_1_3 = lruBit_5_1;
      5'b00110 : _zz__zz_wayToReplace_1_1_3 = lruBit_6_1;
      5'b00111 : _zz__zz_wayToReplace_1_1_3 = lruBit_7_1;
      5'b01000 : _zz__zz_wayToReplace_1_1_3 = lruBit_8_1;
      5'b01001 : _zz__zz_wayToReplace_1_1_3 = lruBit_9_1;
      5'b01010 : _zz__zz_wayToReplace_1_1_3 = lruBit_10_1;
      5'b01011 : _zz__zz_wayToReplace_1_1_3 = lruBit_11_1;
      5'b01100 : _zz__zz_wayToReplace_1_1_3 = lruBit_12_1;
      5'b01101 : _zz__zz_wayToReplace_1_1_3 = lruBit_13_1;
      5'b01110 : _zz__zz_wayToReplace_1_1_3 = lruBit_14_1;
      5'b01111 : _zz__zz_wayToReplace_1_1_3 = lruBit_15_1;
      5'b10000 : _zz__zz_wayToReplace_1_1_3 = lruBit_16_1;
      5'b10001 : _zz__zz_wayToReplace_1_1_3 = lruBit_17_1;
      5'b10010 : _zz__zz_wayToReplace_1_1_3 = lruBit_18_1;
      5'b10011 : _zz__zz_wayToReplace_1_1_3 = lruBit_19_1;
      5'b10100 : _zz__zz_wayToReplace_1_1_3 = lruBit_20_1;
      5'b10101 : _zz__zz_wayToReplace_1_1_3 = lruBit_21_1;
      5'b10110 : _zz__zz_wayToReplace_1_1_3 = lruBit_22_1;
      5'b10111 : _zz__zz_wayToReplace_1_1_3 = lruBit_23_1;
      5'b11000 : _zz__zz_wayToReplace_1_1_3 = lruBit_24_1;
      5'b11001 : _zz__zz_wayToReplace_1_1_3 = lruBit_25_1;
      5'b11010 : _zz__zz_wayToReplace_1_1_3 = lruBit_26_1;
      5'b11011 : _zz__zz_wayToReplace_1_1_3 = lruBit_27_1;
      5'b11100 : _zz__zz_wayToReplace_1_1_3 = lruBit_28_1;
      5'b11101 : _zz__zz_wayToReplace_1_1_3 = lruBit_29_1;
      5'b11110 : _zz__zz_wayToReplace_1_1_3 = lruBit_30_1;
      default : _zz__zz_wayToReplace_1_1_3 = lruBit_31_1;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_1_2_2)
      5'b00000 : _zz__zz_wayToReplace_1_2_1 = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace_1_2_1 = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace_1_2_1 = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace_1_2_1 = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace_1_2_1 = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace_1_2_1 = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace_1_2_1 = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace_1_2_1 = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace_1_2_1 = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace_1_2_1 = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace_1_2_1 = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace_1_2_1 = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace_1_2_1 = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace_1_2_1 = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace_1_2_1 = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace_1_2_1 = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace_1_2_1 = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace_1_2_1 = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace_1_2_1 = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace_1_2_1 = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace_1_2_1 = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace_1_2_1 = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace_1_2_1 = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace_1_2_1 = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace_1_2_1 = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace_1_2_1 = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace_1_2_1 = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace_1_2_1 = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace_1_2_1 = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace_1_2_1 = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace_1_2_1 = lruBit_30_0;
      default : _zz__zz_wayToReplace_1_2_1 = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_1_2_4)
      5'b00000 : _zz__zz_wayToReplace_1_2_3 = lruBit_0_2;
      5'b00001 : _zz__zz_wayToReplace_1_2_3 = lruBit_1_2;
      5'b00010 : _zz__zz_wayToReplace_1_2_3 = lruBit_2_2;
      5'b00011 : _zz__zz_wayToReplace_1_2_3 = lruBit_3_2;
      5'b00100 : _zz__zz_wayToReplace_1_2_3 = lruBit_4_2;
      5'b00101 : _zz__zz_wayToReplace_1_2_3 = lruBit_5_2;
      5'b00110 : _zz__zz_wayToReplace_1_2_3 = lruBit_6_2;
      5'b00111 : _zz__zz_wayToReplace_1_2_3 = lruBit_7_2;
      5'b01000 : _zz__zz_wayToReplace_1_2_3 = lruBit_8_2;
      5'b01001 : _zz__zz_wayToReplace_1_2_3 = lruBit_9_2;
      5'b01010 : _zz__zz_wayToReplace_1_2_3 = lruBit_10_2;
      5'b01011 : _zz__zz_wayToReplace_1_2_3 = lruBit_11_2;
      5'b01100 : _zz__zz_wayToReplace_1_2_3 = lruBit_12_2;
      5'b01101 : _zz__zz_wayToReplace_1_2_3 = lruBit_13_2;
      5'b01110 : _zz__zz_wayToReplace_1_2_3 = lruBit_14_2;
      5'b01111 : _zz__zz_wayToReplace_1_2_3 = lruBit_15_2;
      5'b10000 : _zz__zz_wayToReplace_1_2_3 = lruBit_16_2;
      5'b10001 : _zz__zz_wayToReplace_1_2_3 = lruBit_17_2;
      5'b10010 : _zz__zz_wayToReplace_1_2_3 = lruBit_18_2;
      5'b10011 : _zz__zz_wayToReplace_1_2_3 = lruBit_19_2;
      5'b10100 : _zz__zz_wayToReplace_1_2_3 = lruBit_20_2;
      5'b10101 : _zz__zz_wayToReplace_1_2_3 = lruBit_21_2;
      5'b10110 : _zz__zz_wayToReplace_1_2_3 = lruBit_22_2;
      5'b10111 : _zz__zz_wayToReplace_1_2_3 = lruBit_23_2;
      5'b11000 : _zz__zz_wayToReplace_1_2_3 = lruBit_24_2;
      5'b11001 : _zz__zz_wayToReplace_1_2_3 = lruBit_25_2;
      5'b11010 : _zz__zz_wayToReplace_1_2_3 = lruBit_26_2;
      5'b11011 : _zz__zz_wayToReplace_1_2_3 = lruBit_27_2;
      5'b11100 : _zz__zz_wayToReplace_1_2_3 = lruBit_28_2;
      5'b11101 : _zz__zz_wayToReplace_1_2_3 = lruBit_29_2;
      5'b11110 : _zz__zz_wayToReplace_1_2_3 = lruBit_30_2;
      default : _zz__zz_wayToReplace_1_2_3 = lruBit_31_2;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_1_3_2)
      5'b00000 : _zz__zz_wayToReplace_1_3_1 = lruBit_0_0;
      5'b00001 : _zz__zz_wayToReplace_1_3_1 = lruBit_1_0;
      5'b00010 : _zz__zz_wayToReplace_1_3_1 = lruBit_2_0;
      5'b00011 : _zz__zz_wayToReplace_1_3_1 = lruBit_3_0;
      5'b00100 : _zz__zz_wayToReplace_1_3_1 = lruBit_4_0;
      5'b00101 : _zz__zz_wayToReplace_1_3_1 = lruBit_5_0;
      5'b00110 : _zz__zz_wayToReplace_1_3_1 = lruBit_6_0;
      5'b00111 : _zz__zz_wayToReplace_1_3_1 = lruBit_7_0;
      5'b01000 : _zz__zz_wayToReplace_1_3_1 = lruBit_8_0;
      5'b01001 : _zz__zz_wayToReplace_1_3_1 = lruBit_9_0;
      5'b01010 : _zz__zz_wayToReplace_1_3_1 = lruBit_10_0;
      5'b01011 : _zz__zz_wayToReplace_1_3_1 = lruBit_11_0;
      5'b01100 : _zz__zz_wayToReplace_1_3_1 = lruBit_12_0;
      5'b01101 : _zz__zz_wayToReplace_1_3_1 = lruBit_13_0;
      5'b01110 : _zz__zz_wayToReplace_1_3_1 = lruBit_14_0;
      5'b01111 : _zz__zz_wayToReplace_1_3_1 = lruBit_15_0;
      5'b10000 : _zz__zz_wayToReplace_1_3_1 = lruBit_16_0;
      5'b10001 : _zz__zz_wayToReplace_1_3_1 = lruBit_17_0;
      5'b10010 : _zz__zz_wayToReplace_1_3_1 = lruBit_18_0;
      5'b10011 : _zz__zz_wayToReplace_1_3_1 = lruBit_19_0;
      5'b10100 : _zz__zz_wayToReplace_1_3_1 = lruBit_20_0;
      5'b10101 : _zz__zz_wayToReplace_1_3_1 = lruBit_21_0;
      5'b10110 : _zz__zz_wayToReplace_1_3_1 = lruBit_22_0;
      5'b10111 : _zz__zz_wayToReplace_1_3_1 = lruBit_23_0;
      5'b11000 : _zz__zz_wayToReplace_1_3_1 = lruBit_24_0;
      5'b11001 : _zz__zz_wayToReplace_1_3_1 = lruBit_25_0;
      5'b11010 : _zz__zz_wayToReplace_1_3_1 = lruBit_26_0;
      5'b11011 : _zz__zz_wayToReplace_1_3_1 = lruBit_27_0;
      5'b11100 : _zz__zz_wayToReplace_1_3_1 = lruBit_28_0;
      5'b11101 : _zz__zz_wayToReplace_1_3_1 = lruBit_29_0;
      5'b11110 : _zz__zz_wayToReplace_1_3_1 = lruBit_30_0;
      default : _zz__zz_wayToReplace_1_3_1 = lruBit_31_0;
    endcase
  end

  always @(*) begin
    case(_zz__zz_wayToReplace_1_3_4)
      5'b00000 : _zz__zz_wayToReplace_1_3_3 = lruBit_0_2;
      5'b00001 : _zz__zz_wayToReplace_1_3_3 = lruBit_1_2;
      5'b00010 : _zz__zz_wayToReplace_1_3_3 = lruBit_2_2;
      5'b00011 : _zz__zz_wayToReplace_1_3_3 = lruBit_3_2;
      5'b00100 : _zz__zz_wayToReplace_1_3_3 = lruBit_4_2;
      5'b00101 : _zz__zz_wayToReplace_1_3_3 = lruBit_5_2;
      5'b00110 : _zz__zz_wayToReplace_1_3_3 = lruBit_6_2;
      5'b00111 : _zz__zz_wayToReplace_1_3_3 = lruBit_7_2;
      5'b01000 : _zz__zz_wayToReplace_1_3_3 = lruBit_8_2;
      5'b01001 : _zz__zz_wayToReplace_1_3_3 = lruBit_9_2;
      5'b01010 : _zz__zz_wayToReplace_1_3_3 = lruBit_10_2;
      5'b01011 : _zz__zz_wayToReplace_1_3_3 = lruBit_11_2;
      5'b01100 : _zz__zz_wayToReplace_1_3_3 = lruBit_12_2;
      5'b01101 : _zz__zz_wayToReplace_1_3_3 = lruBit_13_2;
      5'b01110 : _zz__zz_wayToReplace_1_3_3 = lruBit_14_2;
      5'b01111 : _zz__zz_wayToReplace_1_3_3 = lruBit_15_2;
      5'b10000 : _zz__zz_wayToReplace_1_3_3 = lruBit_16_2;
      5'b10001 : _zz__zz_wayToReplace_1_3_3 = lruBit_17_2;
      5'b10010 : _zz__zz_wayToReplace_1_3_3 = lruBit_18_2;
      5'b10011 : _zz__zz_wayToReplace_1_3_3 = lruBit_19_2;
      5'b10100 : _zz__zz_wayToReplace_1_3_3 = lruBit_20_2;
      5'b10101 : _zz__zz_wayToReplace_1_3_3 = lruBit_21_2;
      5'b10110 : _zz__zz_wayToReplace_1_3_3 = lruBit_22_2;
      5'b10111 : _zz__zz_wayToReplace_1_3_3 = lruBit_23_2;
      5'b11000 : _zz__zz_wayToReplace_1_3_3 = lruBit_24_2;
      5'b11001 : _zz__zz_wayToReplace_1_3_3 = lruBit_25_2;
      5'b11010 : _zz__zz_wayToReplace_1_3_3 = lruBit_26_2;
      5'b11011 : _zz__zz_wayToReplace_1_3_3 = lruBit_27_2;
      5'b11100 : _zz__zz_wayToReplace_1_3_3 = lruBit_28_2;
      5'b11101 : _zz__zz_wayToReplace_1_3_3 = lruBit_29_2;
      5'b11110 : _zz__zz_wayToReplace_1_3_3 = lruBit_30_2;
      default : _zz__zz_wayToReplace_1_3_3 = lruBit_31_2;
    endcase
  end

  always @(*) begin
    case(_zz_io_output_availMask_3)
      2'b00 : _zz_io_output_availMask_2 = 2'b00;
      2'b01 : _zz_io_output_availMask_2 = 2'b01;
      2'b10 : _zz_io_output_availMask_2 = 2'b01;
      default : _zz_io_output_availMask_2 = 2'b10;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_0_payload_size)
      LSUSizeOp_byte_1 : io_input_0_payload_size_string = "byte_1  ";
      LSUSizeOp_halfword : io_input_0_payload_size_string = "halfword";
      LSUSizeOp_word : io_input_0_payload_size_string = "word    ";
      default : io_input_0_payload_size_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_input_1_payload_size)
      LSUSizeOp_byte_1 : io_input_1_payload_size_string = "byte_1  ";
      LSUSizeOp_halfword : io_input_1_payload_size_string = "halfword";
      LSUSizeOp_word : io_input_1_payload_size_string = "word    ";
      default : io_input_1_payload_size_string = "????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_1_BOOT : fsm_stateReg_string = "BOOT";
      fsm_enumDef_1_idle : fsm_stateReg_string = "idle";
      fsm_enumDef_1_req : fsm_stateReg_string = "req ";
      fsm_enumDef_1_read : fsm_stateReg_string = "read";
      default : fsm_stateReg_string = "????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_1_BOOT : fsm_stateNext_string = "BOOT";
      fsm_enumDef_1_idle : fsm_stateNext_string = "idle";
      fsm_enumDef_1_req : fsm_stateNext_string = "req ";
      fsm_enumDef_1_read : fsm_stateNext_string = "read";
      default : fsm_stateNext_string = "????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_wr_en = 1'b0;
    if(when_StateMachine_l253_1) begin
      if(when_Cache_l180) begin
        if(when_Cache_l182_3) begin
          _zz_wr_en = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    _zz_wr_en_1 = 1'b0;
    if(when_StateMachine_l253_1) begin
      if(when_Cache_l180) begin
        if(when_Cache_l182_2) begin
          _zz_wr_en_1 = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    _zz_wr_en_2 = 1'b0;
    if(when_StateMachine_l253_1) begin
      if(when_Cache_l180) begin
        if(when_Cache_l182_1) begin
          _zz_wr_en_2 = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    _zz_wr_en_3 = 1'b0;
    if(when_StateMachine_l253_1) begin
      if(when_Cache_l180) begin
        if(when_Cache_l182) begin
          _zz_wr_en_3 = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    _zz_wr_en_4 = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_idle : begin
      end
      fsm_enumDef_1_req : begin
      end
      fsm_enumDef_1_read : begin
        if(when_Cache_l198) begin
          if(when_Cache_l200_3) begin
            if(when_Cache_l201_3) begin
              _zz_wr_en_4 = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_wr_en_5 = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_idle : begin
      end
      fsm_enumDef_1_req : begin
      end
      fsm_enumDef_1_read : begin
        if(when_Cache_l198) begin
          if(when_Cache_l200_2) begin
            if(when_Cache_l201_2) begin
              _zz_wr_en_5 = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_wr_en_6 = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_idle : begin
      end
      fsm_enumDef_1_req : begin
      end
      fsm_enumDef_1_read : begin
        if(when_Cache_l198) begin
          if(when_Cache_l200_1) begin
            if(when_Cache_l201_1) begin
              _zz_wr_en_6 = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_wr_en_7 = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_idle : begin
      end
      fsm_enumDef_1_req : begin
      end
      fsm_enumDef_1_read : begin
        if(when_Cache_l198) begin
          if(when_Cache_l200) begin
            if(when_Cache_l201) begin
              _zz_wr_en_7 = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign cacopEn = ((io_ctrl_cacopStoreTag || io_ctrl_cacopIndexInvalidate) || io_ctrl_cacopHitInvalidate);
  always @(*) begin
    stage1Out_thrown_valid = stage1Out_valid;
    if(io_flush) begin
      stage1Out_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    stage1Out_ready = stage1Out_thrown_ready;
    if(io_flush) begin
      stage1Out_ready = 1'b1;
    end
  end

  assign stage1Out_thrown_payload_branchInfo_0_predictPC = stage1Out_payload_branchInfo_0_predictPC;
  assign stage1Out_thrown_payload_branchInfo_0_predictResult = stage1Out_payload_branchInfo_0_predictResult;
  assign stage1Out_thrown_payload_branchInfo_1_predictPC = stage1Out_payload_branchInfo_1_predictPC;
  assign stage1Out_thrown_payload_branchInfo_1_predictResult = stage1Out_payload_branchInfo_1_predictResult;
  assign stage1Out_thrown_payload_exceptionInfo_0_exception = stage1Out_payload_exceptionInfo_0_exception;
  assign stage1Out_thrown_payload_exceptionInfo_0_eCode = stage1Out_payload_exceptionInfo_0_eCode;
  assign stage1Out_thrown_payload_exceptionInfo_0_eSubCode = stage1Out_payload_exceptionInfo_0_eSubCode;
  assign stage1Out_thrown_payload_exceptionInfo_1_exception = stage1Out_payload_exceptionInfo_1_exception;
  assign stage1Out_thrown_payload_exceptionInfo_1_eCode = stage1Out_payload_exceptionInfo_1_eCode;
  assign stage1Out_thrown_payload_exceptionInfo_1_eSubCode = stage1Out_payload_exceptionInfo_1_eSubCode;
  assign stage1Out_thrown_payload_pc_0 = stage1Out_payload_pc_0;
  assign stage1Out_thrown_payload_pc_1 = stage1Out_payload_pc_1;
  assign stage1Out_thrown_payload_valid = stage1Out_payload_valid;
  assign stage1Out_thrown_payload_tlb_hit = stage1Out_payload_tlb_hit;
  assign stage1Out_thrown_payload_tlb_pageInfo_ppn = stage1Out_payload_tlb_pageInfo_ppn;
  assign stage1Out_thrown_payload_tlb_pageInfo_plv = stage1Out_payload_tlb_pageInfo_plv;
  assign stage1Out_thrown_payload_tlb_pageInfo_mat = stage1Out_payload_tlb_pageInfo_mat;
  assign stage1Out_thrown_payload_tlb_pageInfo_d = stage1Out_payload_tlb_pageInfo_d;
  assign stage1Out_thrown_payload_tlb_pageInfo_v = stage1Out_payload_tlb_pageInfo_v;
  assign stage1Out_thrown_payload_wayValid_0 = stage1Out_payload_wayValid_0;
  assign stage1Out_thrown_payload_wayValid_1 = stage1Out_payload_wayValid_1;
  assign stage1Out_thrown_payload_isStoreTag = stage1Out_payload_isStoreTag;
  assign stage1Out_thrown_payload_isIndexInvalidate = stage1Out_payload_isIndexInvalidate;
  assign stage1Out_thrown_payload_isHitInvalidate = stage1Out_payload_isHitInvalidate;
  always @(*) begin
    stage1Out_thrown_ready = stage1Out_thrown_m2sPipe_ready;
    if(when_Stream_l369) begin
      stage1Out_thrown_ready = 1'b1;
    end
  end

  assign when_Stream_l369 = (! stage1Out_thrown_m2sPipe_valid);
  assign stage1Out_thrown_m2sPipe_valid = stage1Out_thrown_rValid;
  assign stage1Out_thrown_m2sPipe_payload_branchInfo_0_predictPC = stage1Out_thrown_rData_branchInfo_0_predictPC;
  assign stage1Out_thrown_m2sPipe_payload_branchInfo_0_predictResult = stage1Out_thrown_rData_branchInfo_0_predictResult;
  assign stage1Out_thrown_m2sPipe_payload_branchInfo_1_predictPC = stage1Out_thrown_rData_branchInfo_1_predictPC;
  assign stage1Out_thrown_m2sPipe_payload_branchInfo_1_predictResult = stage1Out_thrown_rData_branchInfo_1_predictResult;
  assign stage1Out_thrown_m2sPipe_payload_exceptionInfo_0_exception = stage1Out_thrown_rData_exceptionInfo_0_exception;
  assign stage1Out_thrown_m2sPipe_payload_exceptionInfo_0_eCode = stage1Out_thrown_rData_exceptionInfo_0_eCode;
  assign stage1Out_thrown_m2sPipe_payload_exceptionInfo_0_eSubCode = stage1Out_thrown_rData_exceptionInfo_0_eSubCode;
  assign stage1Out_thrown_m2sPipe_payload_exceptionInfo_1_exception = stage1Out_thrown_rData_exceptionInfo_1_exception;
  assign stage1Out_thrown_m2sPipe_payload_exceptionInfo_1_eCode = stage1Out_thrown_rData_exceptionInfo_1_eCode;
  assign stage1Out_thrown_m2sPipe_payload_exceptionInfo_1_eSubCode = stage1Out_thrown_rData_exceptionInfo_1_eSubCode;
  assign stage1Out_thrown_m2sPipe_payload_pc_0 = stage1Out_thrown_rData_pc_0;
  assign stage1Out_thrown_m2sPipe_payload_pc_1 = stage1Out_thrown_rData_pc_1;
  assign stage1Out_thrown_m2sPipe_payload_valid = stage1Out_thrown_rData_valid;
  assign stage1Out_thrown_m2sPipe_payload_tlb_hit = stage1Out_thrown_rData_tlb_hit;
  assign stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_ppn = stage1Out_thrown_rData_tlb_pageInfo_ppn;
  assign stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_plv = stage1Out_thrown_rData_tlb_pageInfo_plv;
  assign stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_mat = stage1Out_thrown_rData_tlb_pageInfo_mat;
  assign stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_d = stage1Out_thrown_rData_tlb_pageInfo_d;
  assign stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_v = stage1Out_thrown_rData_tlb_pageInfo_v;
  assign stage1Out_thrown_m2sPipe_payload_wayValid_0 = stage1Out_thrown_rData_wayValid_0;
  assign stage1Out_thrown_m2sPipe_payload_wayValid_1 = stage1Out_thrown_rData_wayValid_1;
  assign stage1Out_thrown_m2sPipe_payload_isStoreTag = stage1Out_thrown_rData_isStoreTag;
  assign stage1Out_thrown_m2sPipe_payload_isIndexInvalidate = stage1Out_thrown_rData_isIndexInvalidate;
  assign stage1Out_thrown_m2sPipe_payload_isHitInvalidate = stage1Out_thrown_rData_isHitInvalidate;
  assign stage2In_valid = stage1Out_thrown_m2sPipe_valid;
  assign stage1Out_thrown_m2sPipe_ready = stage2In_ready;
  assign stage2In_payload_branchInfo_0_predictPC = stage1Out_thrown_m2sPipe_payload_branchInfo_0_predictPC;
  assign stage2In_payload_branchInfo_0_predictResult = stage1Out_thrown_m2sPipe_payload_branchInfo_0_predictResult;
  assign stage2In_payload_branchInfo_1_predictPC = stage1Out_thrown_m2sPipe_payload_branchInfo_1_predictPC;
  assign stage2In_payload_branchInfo_1_predictResult = stage1Out_thrown_m2sPipe_payload_branchInfo_1_predictResult;
  assign stage2In_payload_exceptionInfo_0_exception = stage1Out_thrown_m2sPipe_payload_exceptionInfo_0_exception;
  assign stage2In_payload_exceptionInfo_0_eCode = stage1Out_thrown_m2sPipe_payload_exceptionInfo_0_eCode;
  assign stage2In_payload_exceptionInfo_0_eSubCode = stage1Out_thrown_m2sPipe_payload_exceptionInfo_0_eSubCode;
  assign stage2In_payload_exceptionInfo_1_exception = stage1Out_thrown_m2sPipe_payload_exceptionInfo_1_exception;
  assign stage2In_payload_exceptionInfo_1_eCode = stage1Out_thrown_m2sPipe_payload_exceptionInfo_1_eCode;
  assign stage2In_payload_exceptionInfo_1_eSubCode = stage1Out_thrown_m2sPipe_payload_exceptionInfo_1_eSubCode;
  assign stage2In_payload_pc_0 = stage1Out_thrown_m2sPipe_payload_pc_0;
  assign stage2In_payload_pc_1 = stage1Out_thrown_m2sPipe_payload_pc_1;
  assign stage2In_payload_valid = stage1Out_thrown_m2sPipe_payload_valid;
  assign stage2In_payload_tlb_hit = stage1Out_thrown_m2sPipe_payload_tlb_hit;
  assign stage2In_payload_tlb_pageInfo_ppn = stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_ppn;
  assign stage2In_payload_tlb_pageInfo_plv = stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_plv;
  assign stage2In_payload_tlb_pageInfo_mat = stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_mat;
  assign stage2In_payload_tlb_pageInfo_d = stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_d;
  assign stage2In_payload_tlb_pageInfo_v = stage1Out_thrown_m2sPipe_payload_tlb_pageInfo_v;
  assign stage2In_payload_wayValid_0 = stage1Out_thrown_m2sPipe_payload_wayValid_0;
  assign stage2In_payload_wayValid_1 = stage1Out_thrown_m2sPipe_payload_wayValid_1;
  assign stage2In_payload_isStoreTag = stage1Out_thrown_m2sPipe_payload_isStoreTag;
  assign stage2In_payload_isIndexInvalidate = stage1Out_thrown_m2sPipe_payload_isIndexInvalidate;
  assign stage2In_payload_isHitInvalidate = stage1Out_thrown_m2sPipe_payload_isHitInvalidate;
  assign stage1Out_valid = ((|stage1Out_payload_valid) || cacopEn);
  assign io_tlb_virtPageNumber = (io_ctrl_cacopHitInvalidate ? io_ctrl_cacopVA[31 : 12] : io_input_0_payload_address[31 : 12]);
  assign stage1Out_payload_tlb_hit = io_tlb_hit;
  assign stage1Out_payload_tlb_pageInfo_ppn = io_tlb_pageInfo_ppn;
  assign stage1Out_payload_tlb_pageInfo_plv = io_tlb_pageInfo_plv;
  assign stage1Out_payload_tlb_pageInfo_mat = io_tlb_pageInfo_mat;
  assign stage1Out_payload_tlb_pageInfo_d = io_tlb_pageInfo_d;
  assign stage1Out_payload_tlb_pageInfo_v = io_tlb_pageInfo_v;
  assign stage1Out_payload_isStoreTag = io_ctrl_cacopStoreTag;
  assign stage1Out_payload_isIndexInvalidate = io_ctrl_cacopIndexInvalidate;
  assign stage1Out_payload_isHitInvalidate = io_ctrl_cacopHitInvalidate;
  assign stage1Out_fire = (stage1Out_valid && stage1Out_ready);
  assign _zz_io_output_availMask = acceptMask[0];
  assign _zz_io_output_availMask_1 = acceptMask[1];
  always @(*) begin
    stage1Out_payload_wayValid_0[0] = _zz_stage1Out_payload_wayValid_0;
    stage1Out_payload_wayValid_0[1] = _zz_stage1Out_payload_wayValid_0_3;
    stage1Out_payload_wayValid_0[2] = _zz_stage1Out_payload_wayValid_0_6;
    stage1Out_payload_wayValid_0[3] = _zz_stage1Out_payload_wayValid_0_9;
  end

  assign dataRead_0_0 = data_0_rd_data;
  assign tagRead_0_0 = tag_0_rd_data;
  always @(*) begin
    hit_0[0] = ((stage2In_payload_wayValid_0[0] && (tagRead_0_0 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_pc_0[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit_0));
    hit_0[1] = ((stage2In_payload_wayValid_0[1] && (tagRead_0_1 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_pc_0[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit_0_2));
    hit_0[2] = ((stage2In_payload_wayValid_0[2] && (tagRead_0_2 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_pc_0[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit_0_4));
    hit_0[3] = ((stage2In_payload_wayValid_0[3] && (tagRead_0_3 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_pc_0[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit_0_6));
  end

  assign dataRead_0_1 = data_1_rd_data;
  assign tagRead_0_1 = tag_1_rd_data;
  assign dataRead_0_2 = data_2_rd_data;
  assign tagRead_0_2 = tag_2_rd_data;
  assign dataRead_0_3 = data_3_rd_data;
  assign tagRead_0_3 = tag_3_rd_data;
  always @(*) begin
    stage1Out_payload_wayValid_1[0] = _zz_stage1Out_payload_wayValid_1;
    stage1Out_payload_wayValid_1[1] = _zz_stage1Out_payload_wayValid_1_2;
    stage1Out_payload_wayValid_1[2] = _zz_stage1Out_payload_wayValid_1_4;
    stage1Out_payload_wayValid_1[3] = _zz_stage1Out_payload_wayValid_1_6;
  end

  assign dataRead_1_0 = data_0_1_rd_data;
  assign tagRead_1_0 = tag_0_1_rd_data;
  always @(*) begin
    hit_1[0] = ((stage2In_payload_wayValid_1[0] && (tagRead_1_0 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_pc_1[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit_1));
    hit_1[1] = ((stage2In_payload_wayValid_1[1] && (tagRead_1_1 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_pc_1[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit_1_2));
    hit_1[2] = ((stage2In_payload_wayValid_1[2] && (tagRead_1_2 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_pc_1[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit_1_4));
    hit_1[3] = ((stage2In_payload_wayValid_1[3] && (tagRead_1_3 == {stage2In_payload_tlb_pageInfo_ppn,stage2In_payload_pc_1[11 : 11]})) && (stage2In_payload_tlb_pageInfo_mat == _zz_hit_1_6));
  end

  assign dataRead_1_1 = data_1_1_rd_data;
  assign tagRead_1_1 = tag_1_1_rd_data;
  assign dataRead_1_2 = data_2_1_rd_data;
  assign tagRead_1_2 = tag_2_1_rd_data;
  assign dataRead_1_3 = data_3_1_rd_data;
  assign tagRead_1_3 = tag_3_1_rd_data;
  assign fireMask = (io_output_allowMask <<< _zz_fireMask);
  assign stage2In_ready = (((acceptMask | fireMask) == stage2In_payload_valid) || io_flush);
  assign when_Cache_l79 = (! stage2In_payload_tlb_pageInfo_v);
  always @(*) begin
    if(stage2In_payload_tlb_hit) begin
      if(when_Cache_l79) begin
        exceptionInfo2_exception = 1'b1;
      end else begin
        if(when_Cache_l83) begin
          exceptionInfo2_exception = 1'b1;
        end else begin
          exceptionInfo2_exception = 1'b0;
        end
      end
    end else begin
      exceptionInfo2_exception = 1'b1;
    end
  end

  always @(*) begin
    if(stage2In_payload_tlb_hit) begin
      if(when_Cache_l79) begin
        exceptionInfo2_eCode = {4'd0, _zz_exceptionInfo2_eCode};
      end else begin
        if(when_Cache_l83) begin
          exceptionInfo2_eCode = {3'd0, _zz_exceptionInfo2_eCode_1};
        end else begin
          exceptionInfo2_eCode = {3'd0, _zz_exceptionInfo2_eCode_2};
        end
      end
    end else begin
      exceptionInfo2_eCode = 6'h3f;
    end
  end

  always @(*) begin
    if(stage2In_payload_tlb_hit) begin
      if(when_Cache_l79) begin
        exceptionInfo2_eSubCode = 1'b0;
      end else begin
        if(when_Cache_l83) begin
          exceptionInfo2_eSubCode = 1'b0;
        end else begin
          exceptionInfo2_eSubCode = 1'b0;
        end
      end
    end else begin
      exceptionInfo2_eSubCode = 1'b0;
    end
  end

  assign when_Cache_l83 = (stage2In_payload_tlb_pageInfo_plv < _zz_when_Cache_l83);
  assign _zz_missAddr = miss[0];
  assign missAddr = (_zz_missAddr ? stage2In_payload_pc_0 : stage2In_payload_pc_1);
  assign transferAddr = {{stage2In_payload_tlb_pageInfo_ppn,transferIndexOffset},transferBlockOffset};
  always @(*) begin
    miss[0] = (stage2In_payload_valid[0] && (! ((((|hit_0) || io_output_info_0_exceptionInfo_exception) || fetchMask_0) || bufWriteMask[0])));
    miss[1] = (stage2In_payload_valid[1] && (! ((((|hit_1) || io_output_info_1_exceptionInfo_exception) || fetchMask_1) || bufWriteMask[1])));
  end

  always @(*) begin
    sameBlockMask[0] = (io_input_0_valid && (transferAddr[10 : 6] == io_input_0_payload_address[10 : 6]));
    sameBlockMask[1] = (io_input_1_valid && (transferAddr[10 : 6] == io_input_1_payload_address[10 : 6]));
  end

  always @(*) begin
    bufWriteMask[0] = ((io_axi_rvalid && io_axi_rready) && (transferAddr[10 : 0] == stage2In_payload_pc_0[10 : 0]));
    bufWriteMask[1] = ((io_axi_rvalid && io_axi_rready) && (transferAddr[10 : 0] == stage2In_payload_pc_1[10 : 0]));
  end

  assign stall = (io_ctrl_stall || ((|sameBlockMask) && refilling));
  assign when_Cache_l131 = (fireMask[0] && (stage2In_payload_tlb_pageInfo_mat == _zz_when_Cache_l131));
  assign when_Cache_l311 = ((|wayOfReplace_0[3 : 0]) || (|hit_0[3 : 0]));
  assign _zz_1 = ({31'd0,1'b1} <<< stage2In_payload_pc_0[10 : 6]);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = _zz_1[4];
  assign _zz_7 = _zz_1[5];
  assign _zz_8 = _zz_1[6];
  assign _zz_9 = _zz_1[7];
  assign _zz_10 = _zz_1[8];
  assign _zz_11 = _zz_1[9];
  assign _zz_12 = _zz_1[10];
  assign _zz_13 = _zz_1[11];
  assign _zz_14 = _zz_1[12];
  assign _zz_15 = _zz_1[13];
  assign _zz_16 = _zz_1[14];
  assign _zz_17 = _zz_1[15];
  assign _zz_18 = _zz_1[16];
  assign _zz_19 = _zz_1[17];
  assign _zz_20 = _zz_1[18];
  assign _zz_21 = _zz_1[19];
  assign _zz_22 = _zz_1[20];
  assign _zz_23 = _zz_1[21];
  assign _zz_24 = _zz_1[22];
  assign _zz_25 = _zz_1[23];
  assign _zz_26 = _zz_1[24];
  assign _zz_27 = _zz_1[25];
  assign _zz_28 = _zz_1[26];
  assign _zz_29 = _zz_1[27];
  assign _zz_30 = _zz_1[28];
  assign _zz_31 = _zz_1[29];
  assign _zz_32 = _zz_1[30];
  assign _zz_33 = _zz_1[31];
  assign _zz_lruBit_0_0 = ((|wayOfReplace_0[3 : 2]) || (|hit_0[3 : 2]));
  assign when_Cache_l311_1 = ((|wayOfReplace_0[1 : 0]) || (|hit_0[1 : 0]));
  assign _zz_lruBit_0_1 = ((|wayOfReplace_0[1 : 1]) || (|hit_0[1 : 1]));
  assign when_Cache_l311_2 = ((|wayOfReplace_0[3 : 2]) || (|hit_0[3 : 2]));
  assign _zz_lruBit_0_2 = ((|wayOfReplace_0[3 : 3]) || (|hit_0[3 : 3]));
  assign when_Cache_l131_1 = (fireMask[1] && (stage2In_payload_tlb_pageInfo_mat == _zz_when_Cache_l131_1_1));
  assign when_Cache_l311_3 = ((|wayOfReplace_1[3 : 0]) || (|hit_1[3 : 0]));
  assign _zz_34 = ({31'd0,1'b1} <<< stage2In_payload_pc_1[10 : 6]);
  assign _zz_35 = _zz_34[0];
  assign _zz_36 = _zz_34[1];
  assign _zz_37 = _zz_34[2];
  assign _zz_38 = _zz_34[3];
  assign _zz_39 = _zz_34[4];
  assign _zz_40 = _zz_34[5];
  assign _zz_41 = _zz_34[6];
  assign _zz_42 = _zz_34[7];
  assign _zz_43 = _zz_34[8];
  assign _zz_44 = _zz_34[9];
  assign _zz_45 = _zz_34[10];
  assign _zz_46 = _zz_34[11];
  assign _zz_47 = _zz_34[12];
  assign _zz_48 = _zz_34[13];
  assign _zz_49 = _zz_34[14];
  assign _zz_50 = _zz_34[15];
  assign _zz_51 = _zz_34[16];
  assign _zz_52 = _zz_34[17];
  assign _zz_53 = _zz_34[18];
  assign _zz_54 = _zz_34[19];
  assign _zz_55 = _zz_34[20];
  assign _zz_56 = _zz_34[21];
  assign _zz_57 = _zz_34[22];
  assign _zz_58 = _zz_34[23];
  assign _zz_59 = _zz_34[24];
  assign _zz_60 = _zz_34[25];
  assign _zz_61 = _zz_34[26];
  assign _zz_62 = _zz_34[27];
  assign _zz_63 = _zz_34[28];
  assign _zz_64 = _zz_34[29];
  assign _zz_65 = _zz_34[30];
  assign _zz_66 = _zz_34[31];
  assign _zz_lruBit_0_0_1 = ((|wayOfReplace_1[3 : 2]) || (|hit_1[3 : 2]));
  assign when_Cache_l311_4 = ((|wayOfReplace_1[1 : 0]) || (|hit_1[1 : 0]));
  assign _zz_lruBit_0_1_1 = ((|wayOfReplace_1[1 : 1]) || (|hit_1[1 : 1]));
  assign when_Cache_l311_5 = ((|wayOfReplace_1[3 : 2]) || (|hit_1[3 : 2]));
  assign _zz_lruBit_0_2_1 = ((|wayOfReplace_1[3 : 3]) || (|hit_1[3 : 3]));
  assign io_axi_arid = 4'b0000;
  assign io_axi_araddr = transferAddr;
  assign io_axi_arlen = (transferUncached ? 8'h00 : _zz_io_axi_arlen);
  assign io_axi_arsize = 3'b010;
  assign io_axi_arburst = (transferUncached ? 2'b01 : 2'b10);
  assign io_axi_arlock = 2'b00;
  assign io_axi_arcache = 4'b0000;
  assign io_axi_arprot = 3'b000;
  always @(*) begin
    io_axi_arvalid = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_idle : begin
        io_axi_arvalid = 1'b0;
      end
      fsm_enumDef_1_req : begin
        io_axi_arvalid = 1'b1;
      end
      fsm_enumDef_1_read : begin
        io_axi_arvalid = 1'b0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axi_rready = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_idle : begin
        io_axi_rready = 1'b0;
      end
      fsm_enumDef_1_req : begin
        io_axi_rready = 1'b0;
      end
      fsm_enumDef_1_read : begin
        io_axi_rready = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    refilling = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_idle : begin
        refilling = 1'b0;
      end
      fsm_enumDef_1_req : begin
        refilling = 1'b1;
      end
      fsm_enumDef_1_read : begin
        refilling = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_idle : begin
      end
      fsm_enumDef_1_req : begin
      end
      fsm_enumDef_1_read : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  assign when_Cache_l222 = (|io_input_0_payload_address[1 : 0]);
  always @(*) begin
    if(when_Cache_l222) begin
      exceptionInfo1_0_exception = 1'b1;
    end else begin
      exceptionInfo1_0_exception = 1'b0;
    end
  end

  always @(*) begin
    if(when_Cache_l222) begin
      exceptionInfo1_0_eCode = {2'd0, _zz_exceptionInfo1_0_eCode};
    end else begin
      exceptionInfo1_0_eCode = {2'd0, _zz_exceptionInfo1_0_eCode_1};
    end
  end

  always @(*) begin
    if(when_Cache_l222) begin
      exceptionInfo1_0_eSubCode = 1'b0;
    end else begin
      exceptionInfo1_0_eSubCode = 1'b0;
    end
  end

  always @(*) begin
    allowMask[0] = (io_input_0_payload_address[31 : 11] == io_input_0_payload_address[31 : 11]);
    allowMask[1] = (io_input_1_payload_address[31 : 11] == io_input_0_payload_address[31 : 11]);
  end

  assign io_input_0_ready = (((stage1Out_ready && (! stall)) && (&allowMask[0 : 0])) && (! io_flush));
  assign stage1Out_payload_branchInfo_0_predictPC = io_input_0_payload_branchInfo_predictPC;
  assign stage1Out_payload_branchInfo_0_predictResult = io_input_0_payload_branchInfo_predictResult;
  assign stage1Out_payload_exceptionInfo_0_exception = exceptionInfo1_0_exception;
  assign stage1Out_payload_exceptionInfo_0_eCode = exceptionInfo1_0_eCode;
  assign stage1Out_payload_exceptionInfo_0_eSubCode = exceptionInfo1_0_eSubCode;
  assign stage1Out_payload_pc_0 = (cacopEn ? io_ctrl_cacopVA : io_input_0_payload_address);
  assign io_input_0_fire = (io_input_0_valid && io_input_0_ready);
  always @(*) begin
    stage1Out_payload_valid[0] = io_input_0_fire;
    stage1Out_payload_valid[1] = (io_input_1_fire && (io_input_1_payload_address[31 : 11] == io_input_0_payload_address[31 : 11]));
  end

  always @(*) begin
    availMask[0] = (stage2In_payload_valid[0] && (((((|hit_0) || io_output_info_0_exceptionInfo_exception) || acceptMask[0]) || fetchMask_0) || bufWriteMask[0]));
    availMask[1] = (stage2In_payload_valid[1] && (((((|hit_1) || io_output_info_1_exceptionInfo_exception) || acceptMask[1]) || fetchMask_1) || bufWriteMask[1]));
  end

  always @(*) begin
    portAvail[0] = (&availMask[0 : 0]);
    portAvail[1] = (&availMask[1 : 0]);
  end

  assign _zz_portData_0_inst = hit_0[3];
  assign _zz_portData_0_inst_1 = (hit_0[1] || _zz_portData_0_inst);
  assign _zz_portData_0_inst_2 = (hit_0[2] || _zz_portData_0_inst);
  assign portData_0_inst = (((fetchMask_0 || miss[0]) || bufWriteMask[0]) ? (bufWriteMask[0] ? io_axi_rdata : missBuffer_0) : _zz_portData_0_inst_3);
  assign portData_0_branchInfo_predictPC = stage2In_payload_branchInfo_0_predictPC;
  assign portData_0_branchInfo_predictResult = stage2In_payload_branchInfo_0_predictResult;
  assign portData_0_exceptionInfo_exception = (stage2In_payload_exceptionInfo_0_exception ? exceptionInfo2_exception : stage2In_payload_exceptionInfo_0_exception);
  assign portData_0_exceptionInfo_eCode = (stage2In_payload_exceptionInfo_0_exception ? exceptionInfo2_eCode : stage2In_payload_exceptionInfo_0_eCode);
  assign portData_0_exceptionInfo_eSubCode = (stage2In_payload_exceptionInfo_0_exception ? exceptionInfo2_eSubCode : stage2In_payload_exceptionInfo_0_eSubCode);
  assign portData_0_pc = stage2In_payload_pc_0;
  assign when_Cache_l255 = bufWriteMask[0];
  assign _zz_io_output_info_0_inst = _zz__zz_io_output_info_0_inst[0:0];
  assign io_output_info_0_inst = _zz_io_output_info_0_inst_1;
  assign io_output_info_0_branchInfo_predictPC = _zz_io_output_info_0_branchInfo_predictPC;
  assign io_output_info_0_branchInfo_predictResult = _zz_io_output_info_0_branchInfo_predictResult;
  assign io_output_info_0_exceptionInfo_exception = _zz_io_output_info_0_exceptionInfo_exception;
  assign io_output_info_0_exceptionInfo_eCode = _zz_io_output_info_0_exceptionInfo_eCode;
  assign io_output_info_0_exceptionInfo_eSubCode = _zz_io_output_info_0_exceptionInfo_eSubCode;
  assign io_output_info_0_pc = _zz_io_output_info_0_pc;
  always @(*) begin
    hasException[0] = (stage2In_payload_valid[0] && io_output_info_0_exceptionInfo_exception);
    hasException[1] = (stage2In_payload_valid[1] && io_output_info_1_exceptionInfo_exception);
  end

  always @(*) begin
    _zz_wayToReplace_0[0] = (! _zz__zz_wayToReplace_0);
    _zz_wayToReplace_0[1] = (! _zz__zz_wayToReplace_0_2);
  end

  always @(*) begin
    wayToReplace_0[0] = (&_zz_wayToReplace_0);
    wayToReplace_0[1] = (&_zz_wayToReplace_0_1);
    wayToReplace_0[2] = (&_zz_wayToReplace_0_2);
    wayToReplace_0[3] = (&_zz_wayToReplace_0_3);
  end

  always @(*) begin
    _zz_wayToReplace_0_1[0] = (! _zz__zz_wayToReplace_0_1_1);
    _zz_wayToReplace_0_1[1] = _zz__zz_wayToReplace_0_1_3;
  end

  always @(*) begin
    _zz_wayToReplace_0_2[0] = _zz__zz_wayToReplace_0_2_1;
    _zz_wayToReplace_0_2[1] = (! _zz__zz_wayToReplace_0_2_3);
  end

  always @(*) begin
    _zz_wayToReplace_0_3[0] = _zz__zz_wayToReplace_0_3_1;
    _zz_wayToReplace_0_3[1] = _zz__zz_wayToReplace_0_3_3;
  end

  assign when_Cache_l222_1 = (|io_input_1_payload_address[1 : 0]);
  always @(*) begin
    if(when_Cache_l222_1) begin
      exceptionInfo1_1_exception = 1'b1;
    end else begin
      exceptionInfo1_1_exception = 1'b0;
    end
  end

  always @(*) begin
    if(when_Cache_l222_1) begin
      exceptionInfo1_1_eCode = {2'd0, _zz_exceptionInfo1_1_eCode};
    end else begin
      exceptionInfo1_1_eCode = {2'd0, _zz_exceptionInfo1_1_eCode_1};
    end
  end

  always @(*) begin
    if(when_Cache_l222_1) begin
      exceptionInfo1_1_eSubCode = 1'b0;
    end else begin
      exceptionInfo1_1_eSubCode = 1'b0;
    end
  end

  assign io_input_1_ready = (((stage1Out_ready && (! stall)) && (&allowMask[1 : 0])) && (! io_flush));
  assign stage1Out_payload_branchInfo_1_predictPC = io_input_1_payload_branchInfo_predictPC;
  assign stage1Out_payload_branchInfo_1_predictResult = io_input_1_payload_branchInfo_predictResult;
  assign stage1Out_payload_exceptionInfo_1_exception = exceptionInfo1_1_exception;
  assign stage1Out_payload_exceptionInfo_1_eCode = exceptionInfo1_1_eCode;
  assign stage1Out_payload_exceptionInfo_1_eSubCode = exceptionInfo1_1_eSubCode;
  assign stage1Out_payload_pc_1 = io_input_1_payload_address;
  assign io_input_1_fire = (io_input_1_valid && io_input_1_ready);
  assign _zz_portData_1_inst = hit_1[3];
  assign _zz_portData_1_inst_1 = (hit_1[1] || _zz_portData_1_inst);
  assign _zz_portData_1_inst_2 = (hit_1[2] || _zz_portData_1_inst);
  assign portData_1_inst = (((fetchMask_1 || miss[1]) || bufWriteMask[1]) ? (bufWriteMask[1] ? io_axi_rdata : missBuffer_1) : _zz_portData_1_inst_3);
  assign portData_1_branchInfo_predictPC = stage2In_payload_branchInfo_1_predictPC;
  assign portData_1_branchInfo_predictResult = stage2In_payload_branchInfo_1_predictResult;
  assign portData_1_exceptionInfo_exception = (stage2In_payload_exceptionInfo_1_exception ? exceptionInfo2_exception : stage2In_payload_exceptionInfo_1_exception);
  assign portData_1_exceptionInfo_eCode = (stage2In_payload_exceptionInfo_1_exception ? exceptionInfo2_eCode : stage2In_payload_exceptionInfo_1_eCode);
  assign portData_1_exceptionInfo_eSubCode = (stage2In_payload_exceptionInfo_1_exception ? exceptionInfo2_eSubCode : stage2In_payload_exceptionInfo_1_eSubCode);
  assign portData_1_pc = stage2In_payload_pc_1;
  assign when_Cache_l255_1 = bufWriteMask[1];
  assign _zz_io_output_info_1_inst = _zz__zz_io_output_info_1_inst[0:0];
  assign io_output_info_1_inst = _zz_io_output_info_1_inst_1;
  assign io_output_info_1_branchInfo_predictPC = _zz_io_output_info_1_branchInfo_predictPC;
  assign io_output_info_1_branchInfo_predictResult = _zz_io_output_info_1_branchInfo_predictResult;
  assign io_output_info_1_exceptionInfo_exception = _zz_io_output_info_1_exceptionInfo_exception;
  assign io_output_info_1_exceptionInfo_eCode = _zz_io_output_info_1_exceptionInfo_eCode;
  assign io_output_info_1_exceptionInfo_eSubCode = _zz_io_output_info_1_exceptionInfo_eSubCode;
  assign io_output_info_1_pc = _zz_io_output_info_1_pc;
  always @(*) begin
    _zz_wayToReplace_1[0] = (! _zz__zz_wayToReplace_1);
    _zz_wayToReplace_1[1] = (! _zz__zz_wayToReplace_1_2);
  end

  always @(*) begin
    wayToReplace_1[0] = (&_zz_wayToReplace_1);
    wayToReplace_1[1] = (&_zz_wayToReplace_1_1);
    wayToReplace_1[2] = (&_zz_wayToReplace_1_2);
    wayToReplace_1[3] = (&_zz_wayToReplace_1_3);
  end

  always @(*) begin
    _zz_wayToReplace_1_1[0] = (! _zz__zz_wayToReplace_1_1_1);
    _zz_wayToReplace_1_1[1] = _zz__zz_wayToReplace_1_1_3;
  end

  always @(*) begin
    _zz_wayToReplace_1_2[0] = _zz__zz_wayToReplace_1_2_1;
    _zz_wayToReplace_1_2[1] = (! _zz__zz_wayToReplace_1_2_3);
  end

  always @(*) begin
    _zz_wayToReplace_1_3[0] = _zz__zz_wayToReplace_1_3_1;
    _zz_wayToReplace_1_3[1] = _zz__zz_wayToReplace_1_3_3;
  end

  assign io_output_availMask = (portAvail >>> _zz_io_output_availMask_2);
  assign io_badv_vaddr = (hasException[0] ? stage2In_payload_pc_0 : stage2In_payload_pc_1);
  assign io_badv_wen = (|hasException);
  assign io_ctrl_busy = ((refilling || ((|miss) && stage2In_valid)) || (stage2In_valid && ((stage2In_payload_isHitInvalidate || stage2In_payload_isIndexInvalidate) || stage2In_payload_isStoreTag)));
  assign cacopIdx = stage2In_payload_pc_0[10 : 6];
  assign cacopWay = (stage2In_payload_isHitInvalidate ? hit_0 : _zz_cacopWay);
  assign when_Cache_l283 = (stage2In_valid && ((stage2In_payload_isHitInvalidate || stage2In_payload_isIndexInvalidate) || stage2In_payload_isStoreTag));
  assign when_Cache_l285 = cacopWay[0];
  assign _zz_67 = ({31'd0,1'b1} <<< cacopIdx);
  assign when_Cache_l285_1 = cacopWay[1];
  assign _zz_68 = ({31'd0,1'b1} <<< cacopIdx);
  assign when_Cache_l285_2 = cacopWay[2];
  assign _zz_69 = ({31'd0,1'b1} <<< cacopIdx);
  assign when_Cache_l285_3 = cacopWay[3];
  assign _zz_70 = ({31'd0,1'b1} <<< cacopIdx);
  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_enumDef_1_idle : begin
        if(when_Cache_l158) begin
          fsm_stateNext = fsm_enumDef_1_req;
        end
      end
      fsm_enumDef_1_req : begin
        if(when_Cache_l174) begin
          fsm_stateNext = fsm_enumDef_1_read;
        end
      end
      fsm_enumDef_1_read : begin
        if(when_Cache_l209) begin
          if(when_Cache_l210) begin
            fsm_stateNext = fsm_enumDef_1_req;
          end else begin
            fsm_stateNext = fsm_enumDef_1_idle;
          end
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_enumDef_1_idle;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_1_BOOT;
    end
  end

  assign when_Cache_l158 = (((|miss) && stage2In_valid) && (! io_flush));
  assign when_Cache_l174 = (io_axi_arvalid && io_axi_arready);
  assign when_Cache_l198 = (stage2In_payload_tlb_pageInfo_mat == _zz_when_Cache_l198);
  assign when_Cache_l200 = (io_axi_rvalid && io_axi_rready);
  assign when_Cache_l201 = replacingWay[0];
  assign _zz_wr_addr = transferAddr[10 : 2];
  assign _zz_wr_data = io_axi_rdata;
  assign when_Cache_l200_1 = (io_axi_rvalid && io_axi_rready);
  assign when_Cache_l201_1 = replacingWay[1];
  assign _zz_wr_addr_1 = transferAddr[10 : 2];
  assign _zz_wr_data_1 = io_axi_rdata;
  assign when_Cache_l200_2 = (io_axi_rvalid && io_axi_rready);
  assign when_Cache_l201_2 = replacingWay[2];
  assign _zz_wr_addr_2 = transferAddr[10 : 2];
  assign _zz_wr_data_2 = io_axi_rdata;
  assign when_Cache_l200_3 = (io_axi_rvalid && io_axi_rready);
  assign when_Cache_l201_3 = replacingWay[3];
  assign _zz_wr_addr_3 = transferAddr[10 : 2];
  assign _zz_wr_data_3 = io_axi_rdata;
  assign when_Cache_l209 = (io_axi_rlast && (io_axi_rvalid && io_axi_rready));
  assign when_Cache_l210 = (((|miss) && stage2In_valid) && (! io_flush));
  assign when_StateMachine_l253 = ((! (fsm_stateReg == fsm_enumDef_1_req)) && (fsm_stateNext == fsm_enumDef_1_req));
  assign when_StateMachine_l253_1 = ((! (fsm_stateReg == fsm_enumDef_1_read)) && (fsm_stateNext == fsm_enumDef_1_read));
  assign when_Cache_l180 = (stage2In_payload_tlb_pageInfo_mat == _zz_when_Cache_l180);
  assign when_Cache_l182 = replacingWay[0];
  assign _zz_wr_addr_4 = transferAddr[10 : 6];
  assign _zz_wr_data_4 = {stage2In_payload_tlb_pageInfo_ppn,transferAddr[11 : 11]};
  assign _zz_71 = ({31'd0,1'b1} <<< transferAddr[10 : 6]);
  assign when_Cache_l182_1 = replacingWay[1];
  assign _zz_wr_addr_5 = transferAddr[10 : 6];
  assign _zz_wr_data_5 = {stage2In_payload_tlb_pageInfo_ppn,transferAddr[11 : 11]};
  assign _zz_72 = ({31'd0,1'b1} <<< transferAddr[10 : 6]);
  assign when_Cache_l182_2 = replacingWay[2];
  assign _zz_wr_addr_6 = transferAddr[10 : 6];
  assign _zz_wr_data_6 = {stage2In_payload_tlb_pageInfo_ppn,transferAddr[11 : 11]};
  assign _zz_73 = ({31'd0,1'b1} <<< transferAddr[10 : 6]);
  assign when_Cache_l182_3 = replacingWay[3];
  assign _zz_wr_addr_7 = transferAddr[10 : 6];
  assign _zz_wr_data_7 = {stage2In_payload_tlb_pageInfo_ppn,transferAddr[11 : 11]};
  assign _zz_74 = ({31'd0,1'b1} <<< transferAddr[10 : 6]);
  assign when_Cache_l188 = (transferAddr[10 : 6] == stage2In_payload_pc_0[10 : 6]);
  assign when_Cache_l188_1 = (transferAddr[10 : 6] == stage2In_payload_pc_1[10 : 6]);
  assign data_0_wr_en = (_zz_wr_en_7 && 1'b1);
  assign data_0_wr_mask = 1'b1;
  assign data_0_rd_en = (stage1Out_fire && 1'b1);
  assign data_0_rd_addr = _zz_rd_addr[10 : 2];
  assign data_0_1_wr_en = (_zz_wr_en_7 && 1'b1);
  assign data_0_1_wr_mask = 1'b1;
  assign data_0_1_rd_en = (stage1Out_fire && 1'b1);
  assign data_0_1_rd_addr = io_input_1_payload_address[10 : 2];
  assign data_1_wr_en = (_zz_wr_en_6 && 1'b1);
  assign data_1_wr_mask = 1'b1;
  assign data_1_rd_en = (stage1Out_fire && 1'b1);
  assign data_1_rd_addr = _zz_rd_addr_1[10 : 2];
  assign data_1_1_wr_en = (_zz_wr_en_6 && 1'b1);
  assign data_1_1_wr_mask = 1'b1;
  assign data_1_1_rd_en = (stage1Out_fire && 1'b1);
  assign data_1_1_rd_addr = io_input_1_payload_address[10 : 2];
  assign data_2_wr_en = (_zz_wr_en_5 && 1'b1);
  assign data_2_wr_mask = 1'b1;
  assign data_2_rd_en = (stage1Out_fire && 1'b1);
  assign data_2_rd_addr = _zz_rd_addr_2[10 : 2];
  assign data_2_1_wr_en = (_zz_wr_en_5 && 1'b1);
  assign data_2_1_wr_mask = 1'b1;
  assign data_2_1_rd_en = (stage1Out_fire && 1'b1);
  assign data_2_1_rd_addr = io_input_1_payload_address[10 : 2];
  assign data_3_wr_en = (_zz_wr_en_4 && 1'b1);
  assign data_3_wr_mask = 1'b1;
  assign data_3_rd_en = (stage1Out_fire && 1'b1);
  assign data_3_rd_addr = _zz_rd_addr_3[10 : 2];
  assign data_3_1_wr_en = (_zz_wr_en_4 && 1'b1);
  assign data_3_1_wr_mask = 1'b1;
  assign data_3_1_rd_en = (stage1Out_fire && 1'b1);
  assign data_3_1_rd_addr = io_input_1_payload_address[10 : 2];
  assign tag_0_wr_en = (_zz_wr_en_3 && 1'b1);
  assign tag_0_wr_mask = 1'b1;
  assign tag_0_rd_en = (stage1Out_fire && 1'b1);
  assign tag_0_rd_addr = _zz_rd_addr_4[10 : 6];
  assign tag_0_1_wr_en = (_zz_wr_en_3 && 1'b1);
  assign tag_0_1_wr_mask = 1'b1;
  assign tag_0_1_rd_en = (stage1Out_fire && 1'b1);
  assign tag_0_1_rd_addr = io_input_1_payload_address[10 : 6];
  assign tag_1_wr_en = (_zz_wr_en_2 && 1'b1);
  assign tag_1_wr_mask = 1'b1;
  assign tag_1_rd_en = (stage1Out_fire && 1'b1);
  assign tag_1_rd_addr = _zz_rd_addr_5[10 : 6];
  assign tag_1_1_wr_en = (_zz_wr_en_2 && 1'b1);
  assign tag_1_1_wr_mask = 1'b1;
  assign tag_1_1_rd_en = (stage1Out_fire && 1'b1);
  assign tag_1_1_rd_addr = io_input_1_payload_address[10 : 6];
  assign tag_2_wr_en = (_zz_wr_en_1 && 1'b1);
  assign tag_2_wr_mask = 1'b1;
  assign tag_2_rd_en = (stage1Out_fire && 1'b1);
  assign tag_2_rd_addr = _zz_rd_addr_6[10 : 6];
  assign tag_2_1_wr_en = (_zz_wr_en_1 && 1'b1);
  assign tag_2_1_wr_mask = 1'b1;
  assign tag_2_1_rd_en = (stage1Out_fire && 1'b1);
  assign tag_2_1_rd_addr = io_input_1_payload_address[10 : 6];
  assign tag_3_wr_en = (_zz_wr_en && 1'b1);
  assign tag_3_wr_mask = 1'b1;
  assign tag_3_rd_en = (stage1Out_fire && 1'b1);
  assign tag_3_rd_addr = _zz_rd_addr_7[10 : 6];
  assign tag_3_1_wr_en = (_zz_wr_en && 1'b1);
  assign tag_3_1_wr_mask = 1'b1;
  assign tag_3_1_rd_en = (stage1Out_fire && 1'b1);
  assign tag_3_1_rd_addr = io_input_1_payload_address[10 : 6];
  always @(posedge aclk) begin
    if(!aresetn) begin
      valid_0_0 <= 1'b0;
      valid_0_1 <= 1'b0;
      valid_0_2 <= 1'b0;
      valid_0_3 <= 1'b0;
      valid_0_4 <= 1'b0;
      valid_0_5 <= 1'b0;
      valid_0_6 <= 1'b0;
      valid_0_7 <= 1'b0;
      valid_0_8 <= 1'b0;
      valid_0_9 <= 1'b0;
      valid_0_10 <= 1'b0;
      valid_0_11 <= 1'b0;
      valid_0_12 <= 1'b0;
      valid_0_13 <= 1'b0;
      valid_0_14 <= 1'b0;
      valid_0_15 <= 1'b0;
      valid_0_16 <= 1'b0;
      valid_0_17 <= 1'b0;
      valid_0_18 <= 1'b0;
      valid_0_19 <= 1'b0;
      valid_0_20 <= 1'b0;
      valid_0_21 <= 1'b0;
      valid_0_22 <= 1'b0;
      valid_0_23 <= 1'b0;
      valid_0_24 <= 1'b0;
      valid_0_25 <= 1'b0;
      valid_0_26 <= 1'b0;
      valid_0_27 <= 1'b0;
      valid_0_28 <= 1'b0;
      valid_0_29 <= 1'b0;
      valid_0_30 <= 1'b0;
      valid_0_31 <= 1'b0;
      valid_1_0 <= 1'b0;
      valid_1_1 <= 1'b0;
      valid_1_2 <= 1'b0;
      valid_1_3 <= 1'b0;
      valid_1_4 <= 1'b0;
      valid_1_5 <= 1'b0;
      valid_1_6 <= 1'b0;
      valid_1_7 <= 1'b0;
      valid_1_8 <= 1'b0;
      valid_1_9 <= 1'b0;
      valid_1_10 <= 1'b0;
      valid_1_11 <= 1'b0;
      valid_1_12 <= 1'b0;
      valid_1_13 <= 1'b0;
      valid_1_14 <= 1'b0;
      valid_1_15 <= 1'b0;
      valid_1_16 <= 1'b0;
      valid_1_17 <= 1'b0;
      valid_1_18 <= 1'b0;
      valid_1_19 <= 1'b0;
      valid_1_20 <= 1'b0;
      valid_1_21 <= 1'b0;
      valid_1_22 <= 1'b0;
      valid_1_23 <= 1'b0;
      valid_1_24 <= 1'b0;
      valid_1_25 <= 1'b0;
      valid_1_26 <= 1'b0;
      valid_1_27 <= 1'b0;
      valid_1_28 <= 1'b0;
      valid_1_29 <= 1'b0;
      valid_1_30 <= 1'b0;
      valid_1_31 <= 1'b0;
      valid_2_0 <= 1'b0;
      valid_2_1 <= 1'b0;
      valid_2_2 <= 1'b0;
      valid_2_3 <= 1'b0;
      valid_2_4 <= 1'b0;
      valid_2_5 <= 1'b0;
      valid_2_6 <= 1'b0;
      valid_2_7 <= 1'b0;
      valid_2_8 <= 1'b0;
      valid_2_9 <= 1'b0;
      valid_2_10 <= 1'b0;
      valid_2_11 <= 1'b0;
      valid_2_12 <= 1'b0;
      valid_2_13 <= 1'b0;
      valid_2_14 <= 1'b0;
      valid_2_15 <= 1'b0;
      valid_2_16 <= 1'b0;
      valid_2_17 <= 1'b0;
      valid_2_18 <= 1'b0;
      valid_2_19 <= 1'b0;
      valid_2_20 <= 1'b0;
      valid_2_21 <= 1'b0;
      valid_2_22 <= 1'b0;
      valid_2_23 <= 1'b0;
      valid_2_24 <= 1'b0;
      valid_2_25 <= 1'b0;
      valid_2_26 <= 1'b0;
      valid_2_27 <= 1'b0;
      valid_2_28 <= 1'b0;
      valid_2_29 <= 1'b0;
      valid_2_30 <= 1'b0;
      valid_2_31 <= 1'b0;
      valid_3_0 <= 1'b0;
      valid_3_1 <= 1'b0;
      valid_3_2 <= 1'b0;
      valid_3_3 <= 1'b0;
      valid_3_4 <= 1'b0;
      valid_3_5 <= 1'b0;
      valid_3_6 <= 1'b0;
      valid_3_7 <= 1'b0;
      valid_3_8 <= 1'b0;
      valid_3_9 <= 1'b0;
      valid_3_10 <= 1'b0;
      valid_3_11 <= 1'b0;
      valid_3_12 <= 1'b0;
      valid_3_13 <= 1'b0;
      valid_3_14 <= 1'b0;
      valid_3_15 <= 1'b0;
      valid_3_16 <= 1'b0;
      valid_3_17 <= 1'b0;
      valid_3_18 <= 1'b0;
      valid_3_19 <= 1'b0;
      valid_3_20 <= 1'b0;
      valid_3_21 <= 1'b0;
      valid_3_22 <= 1'b0;
      valid_3_23 <= 1'b0;
      valid_3_24 <= 1'b0;
      valid_3_25 <= 1'b0;
      valid_3_26 <= 1'b0;
      valid_3_27 <= 1'b0;
      valid_3_28 <= 1'b0;
      valid_3_29 <= 1'b0;
      valid_3_30 <= 1'b0;
      valid_3_31 <= 1'b0;
      stage1Out_thrown_rValid <= 1'b0;
      acceptMask <= 2'b00;
      lruBit_0_0 <= 1'b0;
      lruBit_0_1 <= 1'b0;
      lruBit_0_2 <= 1'b0;
      lruBit_1_0 <= 1'b0;
      lruBit_1_1 <= 1'b0;
      lruBit_1_2 <= 1'b0;
      lruBit_2_0 <= 1'b0;
      lruBit_2_1 <= 1'b0;
      lruBit_2_2 <= 1'b0;
      lruBit_3_0 <= 1'b0;
      lruBit_3_1 <= 1'b0;
      lruBit_3_2 <= 1'b0;
      lruBit_4_0 <= 1'b0;
      lruBit_4_1 <= 1'b0;
      lruBit_4_2 <= 1'b0;
      lruBit_5_0 <= 1'b0;
      lruBit_5_1 <= 1'b0;
      lruBit_5_2 <= 1'b0;
      lruBit_6_0 <= 1'b0;
      lruBit_6_1 <= 1'b0;
      lruBit_6_2 <= 1'b0;
      lruBit_7_0 <= 1'b0;
      lruBit_7_1 <= 1'b0;
      lruBit_7_2 <= 1'b0;
      lruBit_8_0 <= 1'b0;
      lruBit_8_1 <= 1'b0;
      lruBit_8_2 <= 1'b0;
      lruBit_9_0 <= 1'b0;
      lruBit_9_1 <= 1'b0;
      lruBit_9_2 <= 1'b0;
      lruBit_10_0 <= 1'b0;
      lruBit_10_1 <= 1'b0;
      lruBit_10_2 <= 1'b0;
      lruBit_11_0 <= 1'b0;
      lruBit_11_1 <= 1'b0;
      lruBit_11_2 <= 1'b0;
      lruBit_12_0 <= 1'b0;
      lruBit_12_1 <= 1'b0;
      lruBit_12_2 <= 1'b0;
      lruBit_13_0 <= 1'b0;
      lruBit_13_1 <= 1'b0;
      lruBit_13_2 <= 1'b0;
      lruBit_14_0 <= 1'b0;
      lruBit_14_1 <= 1'b0;
      lruBit_14_2 <= 1'b0;
      lruBit_15_0 <= 1'b0;
      lruBit_15_1 <= 1'b0;
      lruBit_15_2 <= 1'b0;
      lruBit_16_0 <= 1'b0;
      lruBit_16_1 <= 1'b0;
      lruBit_16_2 <= 1'b0;
      lruBit_17_0 <= 1'b0;
      lruBit_17_1 <= 1'b0;
      lruBit_17_2 <= 1'b0;
      lruBit_18_0 <= 1'b0;
      lruBit_18_1 <= 1'b0;
      lruBit_18_2 <= 1'b0;
      lruBit_19_0 <= 1'b0;
      lruBit_19_1 <= 1'b0;
      lruBit_19_2 <= 1'b0;
      lruBit_20_0 <= 1'b0;
      lruBit_20_1 <= 1'b0;
      lruBit_20_2 <= 1'b0;
      lruBit_21_0 <= 1'b0;
      lruBit_21_1 <= 1'b0;
      lruBit_21_2 <= 1'b0;
      lruBit_22_0 <= 1'b0;
      lruBit_22_1 <= 1'b0;
      lruBit_22_2 <= 1'b0;
      lruBit_23_0 <= 1'b0;
      lruBit_23_1 <= 1'b0;
      lruBit_23_2 <= 1'b0;
      lruBit_24_0 <= 1'b0;
      lruBit_24_1 <= 1'b0;
      lruBit_24_2 <= 1'b0;
      lruBit_25_0 <= 1'b0;
      lruBit_25_1 <= 1'b0;
      lruBit_25_2 <= 1'b0;
      lruBit_26_0 <= 1'b0;
      lruBit_26_1 <= 1'b0;
      lruBit_26_2 <= 1'b0;
      lruBit_27_0 <= 1'b0;
      lruBit_27_1 <= 1'b0;
      lruBit_27_2 <= 1'b0;
      lruBit_28_0 <= 1'b0;
      lruBit_28_1 <= 1'b0;
      lruBit_28_2 <= 1'b0;
      lruBit_29_0 <= 1'b0;
      lruBit_29_1 <= 1'b0;
      lruBit_29_2 <= 1'b0;
      lruBit_30_0 <= 1'b0;
      lruBit_30_1 <= 1'b0;
      lruBit_30_2 <= 1'b0;
      lruBit_31_0 <= 1'b0;
      lruBit_31_1 <= 1'b0;
      lruBit_31_2 <= 1'b0;
      fsm_stateReg <= fsm_enumDef_1_BOOT;
    end else begin
      if(stage1Out_thrown_ready) begin
        stage1Out_thrown_rValid <= stage1Out_thrown_valid;
      end
      if(stage1Out_fire) begin
        acceptMask <= 2'b00;
      end else begin
        acceptMask <= (acceptMask | _zz_acceptMask);
      end
      if(when_Cache_l131) begin
        if(when_Cache_l311) begin
          if(_zz_2) begin
            lruBit_0_0 <= _zz_lruBit_0_0;
          end
          if(_zz_3) begin
            lruBit_1_0 <= _zz_lruBit_0_0;
          end
          if(_zz_4) begin
            lruBit_2_0 <= _zz_lruBit_0_0;
          end
          if(_zz_5) begin
            lruBit_3_0 <= _zz_lruBit_0_0;
          end
          if(_zz_6) begin
            lruBit_4_0 <= _zz_lruBit_0_0;
          end
          if(_zz_7) begin
            lruBit_5_0 <= _zz_lruBit_0_0;
          end
          if(_zz_8) begin
            lruBit_6_0 <= _zz_lruBit_0_0;
          end
          if(_zz_9) begin
            lruBit_7_0 <= _zz_lruBit_0_0;
          end
          if(_zz_10) begin
            lruBit_8_0 <= _zz_lruBit_0_0;
          end
          if(_zz_11) begin
            lruBit_9_0 <= _zz_lruBit_0_0;
          end
          if(_zz_12) begin
            lruBit_10_0 <= _zz_lruBit_0_0;
          end
          if(_zz_13) begin
            lruBit_11_0 <= _zz_lruBit_0_0;
          end
          if(_zz_14) begin
            lruBit_12_0 <= _zz_lruBit_0_0;
          end
          if(_zz_15) begin
            lruBit_13_0 <= _zz_lruBit_0_0;
          end
          if(_zz_16) begin
            lruBit_14_0 <= _zz_lruBit_0_0;
          end
          if(_zz_17) begin
            lruBit_15_0 <= _zz_lruBit_0_0;
          end
          if(_zz_18) begin
            lruBit_16_0 <= _zz_lruBit_0_0;
          end
          if(_zz_19) begin
            lruBit_17_0 <= _zz_lruBit_0_0;
          end
          if(_zz_20) begin
            lruBit_18_0 <= _zz_lruBit_0_0;
          end
          if(_zz_21) begin
            lruBit_19_0 <= _zz_lruBit_0_0;
          end
          if(_zz_22) begin
            lruBit_20_0 <= _zz_lruBit_0_0;
          end
          if(_zz_23) begin
            lruBit_21_0 <= _zz_lruBit_0_0;
          end
          if(_zz_24) begin
            lruBit_22_0 <= _zz_lruBit_0_0;
          end
          if(_zz_25) begin
            lruBit_23_0 <= _zz_lruBit_0_0;
          end
          if(_zz_26) begin
            lruBit_24_0 <= _zz_lruBit_0_0;
          end
          if(_zz_27) begin
            lruBit_25_0 <= _zz_lruBit_0_0;
          end
          if(_zz_28) begin
            lruBit_26_0 <= _zz_lruBit_0_0;
          end
          if(_zz_29) begin
            lruBit_27_0 <= _zz_lruBit_0_0;
          end
          if(_zz_30) begin
            lruBit_28_0 <= _zz_lruBit_0_0;
          end
          if(_zz_31) begin
            lruBit_29_0 <= _zz_lruBit_0_0;
          end
          if(_zz_32) begin
            lruBit_30_0 <= _zz_lruBit_0_0;
          end
          if(_zz_33) begin
            lruBit_31_0 <= _zz_lruBit_0_0;
          end
        end
        if(when_Cache_l311_1) begin
          if(_zz_2) begin
            lruBit_0_1 <= _zz_lruBit_0_1;
          end
          if(_zz_3) begin
            lruBit_1_1 <= _zz_lruBit_0_1;
          end
          if(_zz_4) begin
            lruBit_2_1 <= _zz_lruBit_0_1;
          end
          if(_zz_5) begin
            lruBit_3_1 <= _zz_lruBit_0_1;
          end
          if(_zz_6) begin
            lruBit_4_1 <= _zz_lruBit_0_1;
          end
          if(_zz_7) begin
            lruBit_5_1 <= _zz_lruBit_0_1;
          end
          if(_zz_8) begin
            lruBit_6_1 <= _zz_lruBit_0_1;
          end
          if(_zz_9) begin
            lruBit_7_1 <= _zz_lruBit_0_1;
          end
          if(_zz_10) begin
            lruBit_8_1 <= _zz_lruBit_0_1;
          end
          if(_zz_11) begin
            lruBit_9_1 <= _zz_lruBit_0_1;
          end
          if(_zz_12) begin
            lruBit_10_1 <= _zz_lruBit_0_1;
          end
          if(_zz_13) begin
            lruBit_11_1 <= _zz_lruBit_0_1;
          end
          if(_zz_14) begin
            lruBit_12_1 <= _zz_lruBit_0_1;
          end
          if(_zz_15) begin
            lruBit_13_1 <= _zz_lruBit_0_1;
          end
          if(_zz_16) begin
            lruBit_14_1 <= _zz_lruBit_0_1;
          end
          if(_zz_17) begin
            lruBit_15_1 <= _zz_lruBit_0_1;
          end
          if(_zz_18) begin
            lruBit_16_1 <= _zz_lruBit_0_1;
          end
          if(_zz_19) begin
            lruBit_17_1 <= _zz_lruBit_0_1;
          end
          if(_zz_20) begin
            lruBit_18_1 <= _zz_lruBit_0_1;
          end
          if(_zz_21) begin
            lruBit_19_1 <= _zz_lruBit_0_1;
          end
          if(_zz_22) begin
            lruBit_20_1 <= _zz_lruBit_0_1;
          end
          if(_zz_23) begin
            lruBit_21_1 <= _zz_lruBit_0_1;
          end
          if(_zz_24) begin
            lruBit_22_1 <= _zz_lruBit_0_1;
          end
          if(_zz_25) begin
            lruBit_23_1 <= _zz_lruBit_0_1;
          end
          if(_zz_26) begin
            lruBit_24_1 <= _zz_lruBit_0_1;
          end
          if(_zz_27) begin
            lruBit_25_1 <= _zz_lruBit_0_1;
          end
          if(_zz_28) begin
            lruBit_26_1 <= _zz_lruBit_0_1;
          end
          if(_zz_29) begin
            lruBit_27_1 <= _zz_lruBit_0_1;
          end
          if(_zz_30) begin
            lruBit_28_1 <= _zz_lruBit_0_1;
          end
          if(_zz_31) begin
            lruBit_29_1 <= _zz_lruBit_0_1;
          end
          if(_zz_32) begin
            lruBit_30_1 <= _zz_lruBit_0_1;
          end
          if(_zz_33) begin
            lruBit_31_1 <= _zz_lruBit_0_1;
          end
        end
        if(when_Cache_l311_2) begin
          if(_zz_2) begin
            lruBit_0_2 <= _zz_lruBit_0_2;
          end
          if(_zz_3) begin
            lruBit_1_2 <= _zz_lruBit_0_2;
          end
          if(_zz_4) begin
            lruBit_2_2 <= _zz_lruBit_0_2;
          end
          if(_zz_5) begin
            lruBit_3_2 <= _zz_lruBit_0_2;
          end
          if(_zz_6) begin
            lruBit_4_2 <= _zz_lruBit_0_2;
          end
          if(_zz_7) begin
            lruBit_5_2 <= _zz_lruBit_0_2;
          end
          if(_zz_8) begin
            lruBit_6_2 <= _zz_lruBit_0_2;
          end
          if(_zz_9) begin
            lruBit_7_2 <= _zz_lruBit_0_2;
          end
          if(_zz_10) begin
            lruBit_8_2 <= _zz_lruBit_0_2;
          end
          if(_zz_11) begin
            lruBit_9_2 <= _zz_lruBit_0_2;
          end
          if(_zz_12) begin
            lruBit_10_2 <= _zz_lruBit_0_2;
          end
          if(_zz_13) begin
            lruBit_11_2 <= _zz_lruBit_0_2;
          end
          if(_zz_14) begin
            lruBit_12_2 <= _zz_lruBit_0_2;
          end
          if(_zz_15) begin
            lruBit_13_2 <= _zz_lruBit_0_2;
          end
          if(_zz_16) begin
            lruBit_14_2 <= _zz_lruBit_0_2;
          end
          if(_zz_17) begin
            lruBit_15_2 <= _zz_lruBit_0_2;
          end
          if(_zz_18) begin
            lruBit_16_2 <= _zz_lruBit_0_2;
          end
          if(_zz_19) begin
            lruBit_17_2 <= _zz_lruBit_0_2;
          end
          if(_zz_20) begin
            lruBit_18_2 <= _zz_lruBit_0_2;
          end
          if(_zz_21) begin
            lruBit_19_2 <= _zz_lruBit_0_2;
          end
          if(_zz_22) begin
            lruBit_20_2 <= _zz_lruBit_0_2;
          end
          if(_zz_23) begin
            lruBit_21_2 <= _zz_lruBit_0_2;
          end
          if(_zz_24) begin
            lruBit_22_2 <= _zz_lruBit_0_2;
          end
          if(_zz_25) begin
            lruBit_23_2 <= _zz_lruBit_0_2;
          end
          if(_zz_26) begin
            lruBit_24_2 <= _zz_lruBit_0_2;
          end
          if(_zz_27) begin
            lruBit_25_2 <= _zz_lruBit_0_2;
          end
          if(_zz_28) begin
            lruBit_26_2 <= _zz_lruBit_0_2;
          end
          if(_zz_29) begin
            lruBit_27_2 <= _zz_lruBit_0_2;
          end
          if(_zz_30) begin
            lruBit_28_2 <= _zz_lruBit_0_2;
          end
          if(_zz_31) begin
            lruBit_29_2 <= _zz_lruBit_0_2;
          end
          if(_zz_32) begin
            lruBit_30_2 <= _zz_lruBit_0_2;
          end
          if(_zz_33) begin
            lruBit_31_2 <= _zz_lruBit_0_2;
          end
        end
      end
      if(when_Cache_l131_1) begin
        if(when_Cache_l311_3) begin
          if(_zz_35) begin
            lruBit_0_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_36) begin
            lruBit_1_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_37) begin
            lruBit_2_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_38) begin
            lruBit_3_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_39) begin
            lruBit_4_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_40) begin
            lruBit_5_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_41) begin
            lruBit_6_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_42) begin
            lruBit_7_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_43) begin
            lruBit_8_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_44) begin
            lruBit_9_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_45) begin
            lruBit_10_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_46) begin
            lruBit_11_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_47) begin
            lruBit_12_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_48) begin
            lruBit_13_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_49) begin
            lruBit_14_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_50) begin
            lruBit_15_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_51) begin
            lruBit_16_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_52) begin
            lruBit_17_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_53) begin
            lruBit_18_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_54) begin
            lruBit_19_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_55) begin
            lruBit_20_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_56) begin
            lruBit_21_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_57) begin
            lruBit_22_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_58) begin
            lruBit_23_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_59) begin
            lruBit_24_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_60) begin
            lruBit_25_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_61) begin
            lruBit_26_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_62) begin
            lruBit_27_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_63) begin
            lruBit_28_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_64) begin
            lruBit_29_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_65) begin
            lruBit_30_0 <= _zz_lruBit_0_0_1;
          end
          if(_zz_66) begin
            lruBit_31_0 <= _zz_lruBit_0_0_1;
          end
        end
        if(when_Cache_l311_4) begin
          if(_zz_35) begin
            lruBit_0_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_36) begin
            lruBit_1_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_37) begin
            lruBit_2_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_38) begin
            lruBit_3_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_39) begin
            lruBit_4_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_40) begin
            lruBit_5_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_41) begin
            lruBit_6_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_42) begin
            lruBit_7_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_43) begin
            lruBit_8_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_44) begin
            lruBit_9_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_45) begin
            lruBit_10_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_46) begin
            lruBit_11_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_47) begin
            lruBit_12_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_48) begin
            lruBit_13_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_49) begin
            lruBit_14_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_50) begin
            lruBit_15_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_51) begin
            lruBit_16_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_52) begin
            lruBit_17_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_53) begin
            lruBit_18_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_54) begin
            lruBit_19_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_55) begin
            lruBit_20_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_56) begin
            lruBit_21_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_57) begin
            lruBit_22_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_58) begin
            lruBit_23_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_59) begin
            lruBit_24_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_60) begin
            lruBit_25_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_61) begin
            lruBit_26_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_62) begin
            lruBit_27_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_63) begin
            lruBit_28_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_64) begin
            lruBit_29_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_65) begin
            lruBit_30_1 <= _zz_lruBit_0_1_1;
          end
          if(_zz_66) begin
            lruBit_31_1 <= _zz_lruBit_0_1_1;
          end
        end
        if(when_Cache_l311_5) begin
          if(_zz_35) begin
            lruBit_0_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_36) begin
            lruBit_1_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_37) begin
            lruBit_2_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_38) begin
            lruBit_3_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_39) begin
            lruBit_4_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_40) begin
            lruBit_5_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_41) begin
            lruBit_6_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_42) begin
            lruBit_7_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_43) begin
            lruBit_8_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_44) begin
            lruBit_9_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_45) begin
            lruBit_10_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_46) begin
            lruBit_11_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_47) begin
            lruBit_12_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_48) begin
            lruBit_13_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_49) begin
            lruBit_14_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_50) begin
            lruBit_15_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_51) begin
            lruBit_16_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_52) begin
            lruBit_17_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_53) begin
            lruBit_18_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_54) begin
            lruBit_19_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_55) begin
            lruBit_20_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_56) begin
            lruBit_21_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_57) begin
            lruBit_22_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_58) begin
            lruBit_23_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_59) begin
            lruBit_24_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_60) begin
            lruBit_25_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_61) begin
            lruBit_26_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_62) begin
            lruBit_27_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_63) begin
            lruBit_28_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_64) begin
            lruBit_29_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_65) begin
            lruBit_30_2 <= _zz_lruBit_0_2_1;
          end
          if(_zz_66) begin
            lruBit_31_2 <= _zz_lruBit_0_2_1;
          end
        end
      end
      if(when_Cache_l283) begin
        if(when_Cache_l285) begin
          if(_zz_67[0]) begin
            valid_0_0 <= 1'b0;
          end
          if(_zz_67[1]) begin
            valid_0_1 <= 1'b0;
          end
          if(_zz_67[2]) begin
            valid_0_2 <= 1'b0;
          end
          if(_zz_67[3]) begin
            valid_0_3 <= 1'b0;
          end
          if(_zz_67[4]) begin
            valid_0_4 <= 1'b0;
          end
          if(_zz_67[5]) begin
            valid_0_5 <= 1'b0;
          end
          if(_zz_67[6]) begin
            valid_0_6 <= 1'b0;
          end
          if(_zz_67[7]) begin
            valid_0_7 <= 1'b0;
          end
          if(_zz_67[8]) begin
            valid_0_8 <= 1'b0;
          end
          if(_zz_67[9]) begin
            valid_0_9 <= 1'b0;
          end
          if(_zz_67[10]) begin
            valid_0_10 <= 1'b0;
          end
          if(_zz_67[11]) begin
            valid_0_11 <= 1'b0;
          end
          if(_zz_67[12]) begin
            valid_0_12 <= 1'b0;
          end
          if(_zz_67[13]) begin
            valid_0_13 <= 1'b0;
          end
          if(_zz_67[14]) begin
            valid_0_14 <= 1'b0;
          end
          if(_zz_67[15]) begin
            valid_0_15 <= 1'b0;
          end
          if(_zz_67[16]) begin
            valid_0_16 <= 1'b0;
          end
          if(_zz_67[17]) begin
            valid_0_17 <= 1'b0;
          end
          if(_zz_67[18]) begin
            valid_0_18 <= 1'b0;
          end
          if(_zz_67[19]) begin
            valid_0_19 <= 1'b0;
          end
          if(_zz_67[20]) begin
            valid_0_20 <= 1'b0;
          end
          if(_zz_67[21]) begin
            valid_0_21 <= 1'b0;
          end
          if(_zz_67[22]) begin
            valid_0_22 <= 1'b0;
          end
          if(_zz_67[23]) begin
            valid_0_23 <= 1'b0;
          end
          if(_zz_67[24]) begin
            valid_0_24 <= 1'b0;
          end
          if(_zz_67[25]) begin
            valid_0_25 <= 1'b0;
          end
          if(_zz_67[26]) begin
            valid_0_26 <= 1'b0;
          end
          if(_zz_67[27]) begin
            valid_0_27 <= 1'b0;
          end
          if(_zz_67[28]) begin
            valid_0_28 <= 1'b0;
          end
          if(_zz_67[29]) begin
            valid_0_29 <= 1'b0;
          end
          if(_zz_67[30]) begin
            valid_0_30 <= 1'b0;
          end
          if(_zz_67[31]) begin
            valid_0_31 <= 1'b0;
          end
        end
        if(when_Cache_l285_1) begin
          if(_zz_68[0]) begin
            valid_1_0 <= 1'b0;
          end
          if(_zz_68[1]) begin
            valid_1_1 <= 1'b0;
          end
          if(_zz_68[2]) begin
            valid_1_2 <= 1'b0;
          end
          if(_zz_68[3]) begin
            valid_1_3 <= 1'b0;
          end
          if(_zz_68[4]) begin
            valid_1_4 <= 1'b0;
          end
          if(_zz_68[5]) begin
            valid_1_5 <= 1'b0;
          end
          if(_zz_68[6]) begin
            valid_1_6 <= 1'b0;
          end
          if(_zz_68[7]) begin
            valid_1_7 <= 1'b0;
          end
          if(_zz_68[8]) begin
            valid_1_8 <= 1'b0;
          end
          if(_zz_68[9]) begin
            valid_1_9 <= 1'b0;
          end
          if(_zz_68[10]) begin
            valid_1_10 <= 1'b0;
          end
          if(_zz_68[11]) begin
            valid_1_11 <= 1'b0;
          end
          if(_zz_68[12]) begin
            valid_1_12 <= 1'b0;
          end
          if(_zz_68[13]) begin
            valid_1_13 <= 1'b0;
          end
          if(_zz_68[14]) begin
            valid_1_14 <= 1'b0;
          end
          if(_zz_68[15]) begin
            valid_1_15 <= 1'b0;
          end
          if(_zz_68[16]) begin
            valid_1_16 <= 1'b0;
          end
          if(_zz_68[17]) begin
            valid_1_17 <= 1'b0;
          end
          if(_zz_68[18]) begin
            valid_1_18 <= 1'b0;
          end
          if(_zz_68[19]) begin
            valid_1_19 <= 1'b0;
          end
          if(_zz_68[20]) begin
            valid_1_20 <= 1'b0;
          end
          if(_zz_68[21]) begin
            valid_1_21 <= 1'b0;
          end
          if(_zz_68[22]) begin
            valid_1_22 <= 1'b0;
          end
          if(_zz_68[23]) begin
            valid_1_23 <= 1'b0;
          end
          if(_zz_68[24]) begin
            valid_1_24 <= 1'b0;
          end
          if(_zz_68[25]) begin
            valid_1_25 <= 1'b0;
          end
          if(_zz_68[26]) begin
            valid_1_26 <= 1'b0;
          end
          if(_zz_68[27]) begin
            valid_1_27 <= 1'b0;
          end
          if(_zz_68[28]) begin
            valid_1_28 <= 1'b0;
          end
          if(_zz_68[29]) begin
            valid_1_29 <= 1'b0;
          end
          if(_zz_68[30]) begin
            valid_1_30 <= 1'b0;
          end
          if(_zz_68[31]) begin
            valid_1_31 <= 1'b0;
          end
        end
        if(when_Cache_l285_2) begin
          if(_zz_69[0]) begin
            valid_2_0 <= 1'b0;
          end
          if(_zz_69[1]) begin
            valid_2_1 <= 1'b0;
          end
          if(_zz_69[2]) begin
            valid_2_2 <= 1'b0;
          end
          if(_zz_69[3]) begin
            valid_2_3 <= 1'b0;
          end
          if(_zz_69[4]) begin
            valid_2_4 <= 1'b0;
          end
          if(_zz_69[5]) begin
            valid_2_5 <= 1'b0;
          end
          if(_zz_69[6]) begin
            valid_2_6 <= 1'b0;
          end
          if(_zz_69[7]) begin
            valid_2_7 <= 1'b0;
          end
          if(_zz_69[8]) begin
            valid_2_8 <= 1'b0;
          end
          if(_zz_69[9]) begin
            valid_2_9 <= 1'b0;
          end
          if(_zz_69[10]) begin
            valid_2_10 <= 1'b0;
          end
          if(_zz_69[11]) begin
            valid_2_11 <= 1'b0;
          end
          if(_zz_69[12]) begin
            valid_2_12 <= 1'b0;
          end
          if(_zz_69[13]) begin
            valid_2_13 <= 1'b0;
          end
          if(_zz_69[14]) begin
            valid_2_14 <= 1'b0;
          end
          if(_zz_69[15]) begin
            valid_2_15 <= 1'b0;
          end
          if(_zz_69[16]) begin
            valid_2_16 <= 1'b0;
          end
          if(_zz_69[17]) begin
            valid_2_17 <= 1'b0;
          end
          if(_zz_69[18]) begin
            valid_2_18 <= 1'b0;
          end
          if(_zz_69[19]) begin
            valid_2_19 <= 1'b0;
          end
          if(_zz_69[20]) begin
            valid_2_20 <= 1'b0;
          end
          if(_zz_69[21]) begin
            valid_2_21 <= 1'b0;
          end
          if(_zz_69[22]) begin
            valid_2_22 <= 1'b0;
          end
          if(_zz_69[23]) begin
            valid_2_23 <= 1'b0;
          end
          if(_zz_69[24]) begin
            valid_2_24 <= 1'b0;
          end
          if(_zz_69[25]) begin
            valid_2_25 <= 1'b0;
          end
          if(_zz_69[26]) begin
            valid_2_26 <= 1'b0;
          end
          if(_zz_69[27]) begin
            valid_2_27 <= 1'b0;
          end
          if(_zz_69[28]) begin
            valid_2_28 <= 1'b0;
          end
          if(_zz_69[29]) begin
            valid_2_29 <= 1'b0;
          end
          if(_zz_69[30]) begin
            valid_2_30 <= 1'b0;
          end
          if(_zz_69[31]) begin
            valid_2_31 <= 1'b0;
          end
        end
        if(when_Cache_l285_3) begin
          if(_zz_70[0]) begin
            valid_3_0 <= 1'b0;
          end
          if(_zz_70[1]) begin
            valid_3_1 <= 1'b0;
          end
          if(_zz_70[2]) begin
            valid_3_2 <= 1'b0;
          end
          if(_zz_70[3]) begin
            valid_3_3 <= 1'b0;
          end
          if(_zz_70[4]) begin
            valid_3_4 <= 1'b0;
          end
          if(_zz_70[5]) begin
            valid_3_5 <= 1'b0;
          end
          if(_zz_70[6]) begin
            valid_3_6 <= 1'b0;
          end
          if(_zz_70[7]) begin
            valid_3_7 <= 1'b0;
          end
          if(_zz_70[8]) begin
            valid_3_8 <= 1'b0;
          end
          if(_zz_70[9]) begin
            valid_3_9 <= 1'b0;
          end
          if(_zz_70[10]) begin
            valid_3_10 <= 1'b0;
          end
          if(_zz_70[11]) begin
            valid_3_11 <= 1'b0;
          end
          if(_zz_70[12]) begin
            valid_3_12 <= 1'b0;
          end
          if(_zz_70[13]) begin
            valid_3_13 <= 1'b0;
          end
          if(_zz_70[14]) begin
            valid_3_14 <= 1'b0;
          end
          if(_zz_70[15]) begin
            valid_3_15 <= 1'b0;
          end
          if(_zz_70[16]) begin
            valid_3_16 <= 1'b0;
          end
          if(_zz_70[17]) begin
            valid_3_17 <= 1'b0;
          end
          if(_zz_70[18]) begin
            valid_3_18 <= 1'b0;
          end
          if(_zz_70[19]) begin
            valid_3_19 <= 1'b0;
          end
          if(_zz_70[20]) begin
            valid_3_20 <= 1'b0;
          end
          if(_zz_70[21]) begin
            valid_3_21 <= 1'b0;
          end
          if(_zz_70[22]) begin
            valid_3_22 <= 1'b0;
          end
          if(_zz_70[23]) begin
            valid_3_23 <= 1'b0;
          end
          if(_zz_70[24]) begin
            valid_3_24 <= 1'b0;
          end
          if(_zz_70[25]) begin
            valid_3_25 <= 1'b0;
          end
          if(_zz_70[26]) begin
            valid_3_26 <= 1'b0;
          end
          if(_zz_70[27]) begin
            valid_3_27 <= 1'b0;
          end
          if(_zz_70[28]) begin
            valid_3_28 <= 1'b0;
          end
          if(_zz_70[29]) begin
            valid_3_29 <= 1'b0;
          end
          if(_zz_70[30]) begin
            valid_3_30 <= 1'b0;
          end
          if(_zz_70[31]) begin
            valid_3_31 <= 1'b0;
          end
        end
      end
      fsm_stateReg <= fsm_stateNext;
      if(when_StateMachine_l253_1) begin
        if(when_Cache_l180) begin
          if(when_Cache_l182) begin
            if(_zz_71[0]) begin
              valid_0_0 <= 1'b1;
            end
            if(_zz_71[1]) begin
              valid_0_1 <= 1'b1;
            end
            if(_zz_71[2]) begin
              valid_0_2 <= 1'b1;
            end
            if(_zz_71[3]) begin
              valid_0_3 <= 1'b1;
            end
            if(_zz_71[4]) begin
              valid_0_4 <= 1'b1;
            end
            if(_zz_71[5]) begin
              valid_0_5 <= 1'b1;
            end
            if(_zz_71[6]) begin
              valid_0_6 <= 1'b1;
            end
            if(_zz_71[7]) begin
              valid_0_7 <= 1'b1;
            end
            if(_zz_71[8]) begin
              valid_0_8 <= 1'b1;
            end
            if(_zz_71[9]) begin
              valid_0_9 <= 1'b1;
            end
            if(_zz_71[10]) begin
              valid_0_10 <= 1'b1;
            end
            if(_zz_71[11]) begin
              valid_0_11 <= 1'b1;
            end
            if(_zz_71[12]) begin
              valid_0_12 <= 1'b1;
            end
            if(_zz_71[13]) begin
              valid_0_13 <= 1'b1;
            end
            if(_zz_71[14]) begin
              valid_0_14 <= 1'b1;
            end
            if(_zz_71[15]) begin
              valid_0_15 <= 1'b1;
            end
            if(_zz_71[16]) begin
              valid_0_16 <= 1'b1;
            end
            if(_zz_71[17]) begin
              valid_0_17 <= 1'b1;
            end
            if(_zz_71[18]) begin
              valid_0_18 <= 1'b1;
            end
            if(_zz_71[19]) begin
              valid_0_19 <= 1'b1;
            end
            if(_zz_71[20]) begin
              valid_0_20 <= 1'b1;
            end
            if(_zz_71[21]) begin
              valid_0_21 <= 1'b1;
            end
            if(_zz_71[22]) begin
              valid_0_22 <= 1'b1;
            end
            if(_zz_71[23]) begin
              valid_0_23 <= 1'b1;
            end
            if(_zz_71[24]) begin
              valid_0_24 <= 1'b1;
            end
            if(_zz_71[25]) begin
              valid_0_25 <= 1'b1;
            end
            if(_zz_71[26]) begin
              valid_0_26 <= 1'b1;
            end
            if(_zz_71[27]) begin
              valid_0_27 <= 1'b1;
            end
            if(_zz_71[28]) begin
              valid_0_28 <= 1'b1;
            end
            if(_zz_71[29]) begin
              valid_0_29 <= 1'b1;
            end
            if(_zz_71[30]) begin
              valid_0_30 <= 1'b1;
            end
            if(_zz_71[31]) begin
              valid_0_31 <= 1'b1;
            end
          end
          if(when_Cache_l182_1) begin
            if(_zz_72[0]) begin
              valid_1_0 <= 1'b1;
            end
            if(_zz_72[1]) begin
              valid_1_1 <= 1'b1;
            end
            if(_zz_72[2]) begin
              valid_1_2 <= 1'b1;
            end
            if(_zz_72[3]) begin
              valid_1_3 <= 1'b1;
            end
            if(_zz_72[4]) begin
              valid_1_4 <= 1'b1;
            end
            if(_zz_72[5]) begin
              valid_1_5 <= 1'b1;
            end
            if(_zz_72[6]) begin
              valid_1_6 <= 1'b1;
            end
            if(_zz_72[7]) begin
              valid_1_7 <= 1'b1;
            end
            if(_zz_72[8]) begin
              valid_1_8 <= 1'b1;
            end
            if(_zz_72[9]) begin
              valid_1_9 <= 1'b1;
            end
            if(_zz_72[10]) begin
              valid_1_10 <= 1'b1;
            end
            if(_zz_72[11]) begin
              valid_1_11 <= 1'b1;
            end
            if(_zz_72[12]) begin
              valid_1_12 <= 1'b1;
            end
            if(_zz_72[13]) begin
              valid_1_13 <= 1'b1;
            end
            if(_zz_72[14]) begin
              valid_1_14 <= 1'b1;
            end
            if(_zz_72[15]) begin
              valid_1_15 <= 1'b1;
            end
            if(_zz_72[16]) begin
              valid_1_16 <= 1'b1;
            end
            if(_zz_72[17]) begin
              valid_1_17 <= 1'b1;
            end
            if(_zz_72[18]) begin
              valid_1_18 <= 1'b1;
            end
            if(_zz_72[19]) begin
              valid_1_19 <= 1'b1;
            end
            if(_zz_72[20]) begin
              valid_1_20 <= 1'b1;
            end
            if(_zz_72[21]) begin
              valid_1_21 <= 1'b1;
            end
            if(_zz_72[22]) begin
              valid_1_22 <= 1'b1;
            end
            if(_zz_72[23]) begin
              valid_1_23 <= 1'b1;
            end
            if(_zz_72[24]) begin
              valid_1_24 <= 1'b1;
            end
            if(_zz_72[25]) begin
              valid_1_25 <= 1'b1;
            end
            if(_zz_72[26]) begin
              valid_1_26 <= 1'b1;
            end
            if(_zz_72[27]) begin
              valid_1_27 <= 1'b1;
            end
            if(_zz_72[28]) begin
              valid_1_28 <= 1'b1;
            end
            if(_zz_72[29]) begin
              valid_1_29 <= 1'b1;
            end
            if(_zz_72[30]) begin
              valid_1_30 <= 1'b1;
            end
            if(_zz_72[31]) begin
              valid_1_31 <= 1'b1;
            end
          end
          if(when_Cache_l182_2) begin
            if(_zz_73[0]) begin
              valid_2_0 <= 1'b1;
            end
            if(_zz_73[1]) begin
              valid_2_1 <= 1'b1;
            end
            if(_zz_73[2]) begin
              valid_2_2 <= 1'b1;
            end
            if(_zz_73[3]) begin
              valid_2_3 <= 1'b1;
            end
            if(_zz_73[4]) begin
              valid_2_4 <= 1'b1;
            end
            if(_zz_73[5]) begin
              valid_2_5 <= 1'b1;
            end
            if(_zz_73[6]) begin
              valid_2_6 <= 1'b1;
            end
            if(_zz_73[7]) begin
              valid_2_7 <= 1'b1;
            end
            if(_zz_73[8]) begin
              valid_2_8 <= 1'b1;
            end
            if(_zz_73[9]) begin
              valid_2_9 <= 1'b1;
            end
            if(_zz_73[10]) begin
              valid_2_10 <= 1'b1;
            end
            if(_zz_73[11]) begin
              valid_2_11 <= 1'b1;
            end
            if(_zz_73[12]) begin
              valid_2_12 <= 1'b1;
            end
            if(_zz_73[13]) begin
              valid_2_13 <= 1'b1;
            end
            if(_zz_73[14]) begin
              valid_2_14 <= 1'b1;
            end
            if(_zz_73[15]) begin
              valid_2_15 <= 1'b1;
            end
            if(_zz_73[16]) begin
              valid_2_16 <= 1'b1;
            end
            if(_zz_73[17]) begin
              valid_2_17 <= 1'b1;
            end
            if(_zz_73[18]) begin
              valid_2_18 <= 1'b1;
            end
            if(_zz_73[19]) begin
              valid_2_19 <= 1'b1;
            end
            if(_zz_73[20]) begin
              valid_2_20 <= 1'b1;
            end
            if(_zz_73[21]) begin
              valid_2_21 <= 1'b1;
            end
            if(_zz_73[22]) begin
              valid_2_22 <= 1'b1;
            end
            if(_zz_73[23]) begin
              valid_2_23 <= 1'b1;
            end
            if(_zz_73[24]) begin
              valid_2_24 <= 1'b1;
            end
            if(_zz_73[25]) begin
              valid_2_25 <= 1'b1;
            end
            if(_zz_73[26]) begin
              valid_2_26 <= 1'b1;
            end
            if(_zz_73[27]) begin
              valid_2_27 <= 1'b1;
            end
            if(_zz_73[28]) begin
              valid_2_28 <= 1'b1;
            end
            if(_zz_73[29]) begin
              valid_2_29 <= 1'b1;
            end
            if(_zz_73[30]) begin
              valid_2_30 <= 1'b1;
            end
            if(_zz_73[31]) begin
              valid_2_31 <= 1'b1;
            end
          end
          if(when_Cache_l182_3) begin
            if(_zz_74[0]) begin
              valid_3_0 <= 1'b1;
            end
            if(_zz_74[1]) begin
              valid_3_1 <= 1'b1;
            end
            if(_zz_74[2]) begin
              valid_3_2 <= 1'b1;
            end
            if(_zz_74[3]) begin
              valid_3_3 <= 1'b1;
            end
            if(_zz_74[4]) begin
              valid_3_4 <= 1'b1;
            end
            if(_zz_74[5]) begin
              valid_3_5 <= 1'b1;
            end
            if(_zz_74[6]) begin
              valid_3_6 <= 1'b1;
            end
            if(_zz_74[7]) begin
              valid_3_7 <= 1'b1;
            end
            if(_zz_74[8]) begin
              valid_3_8 <= 1'b1;
            end
            if(_zz_74[9]) begin
              valid_3_9 <= 1'b1;
            end
            if(_zz_74[10]) begin
              valid_3_10 <= 1'b1;
            end
            if(_zz_74[11]) begin
              valid_3_11 <= 1'b1;
            end
            if(_zz_74[12]) begin
              valid_3_12 <= 1'b1;
            end
            if(_zz_74[13]) begin
              valid_3_13 <= 1'b1;
            end
            if(_zz_74[14]) begin
              valid_3_14 <= 1'b1;
            end
            if(_zz_74[15]) begin
              valid_3_15 <= 1'b1;
            end
            if(_zz_74[16]) begin
              valid_3_16 <= 1'b1;
            end
            if(_zz_74[17]) begin
              valid_3_17 <= 1'b1;
            end
            if(_zz_74[18]) begin
              valid_3_18 <= 1'b1;
            end
            if(_zz_74[19]) begin
              valid_3_19 <= 1'b1;
            end
            if(_zz_74[20]) begin
              valid_3_20 <= 1'b1;
            end
            if(_zz_74[21]) begin
              valid_3_21 <= 1'b1;
            end
            if(_zz_74[22]) begin
              valid_3_22 <= 1'b1;
            end
            if(_zz_74[23]) begin
              valid_3_23 <= 1'b1;
            end
            if(_zz_74[24]) begin
              valid_3_24 <= 1'b1;
            end
            if(_zz_74[25]) begin
              valid_3_25 <= 1'b1;
            end
            if(_zz_74[26]) begin
              valid_3_26 <= 1'b1;
            end
            if(_zz_74[27]) begin
              valid_3_27 <= 1'b1;
            end
            if(_zz_74[28]) begin
              valid_3_28 <= 1'b1;
            end
            if(_zz_74[29]) begin
              valid_3_29 <= 1'b1;
            end
            if(_zz_74[30]) begin
              valid_3_30 <= 1'b1;
            end
            if(_zz_74[31]) begin
              valid_3_31 <= 1'b1;
            end
          end
        end
      end
    end
  end

  always @(posedge aclk) begin
    if(stage1Out_thrown_ready) begin
      stage1Out_thrown_rData_branchInfo_0_predictPC <= stage1Out_thrown_payload_branchInfo_0_predictPC;
      stage1Out_thrown_rData_branchInfo_0_predictResult <= stage1Out_thrown_payload_branchInfo_0_predictResult;
      stage1Out_thrown_rData_branchInfo_1_predictPC <= stage1Out_thrown_payload_branchInfo_1_predictPC;
      stage1Out_thrown_rData_branchInfo_1_predictResult <= stage1Out_thrown_payload_branchInfo_1_predictResult;
      stage1Out_thrown_rData_exceptionInfo_0_exception <= stage1Out_thrown_payload_exceptionInfo_0_exception;
      stage1Out_thrown_rData_exceptionInfo_0_eCode <= stage1Out_thrown_payload_exceptionInfo_0_eCode;
      stage1Out_thrown_rData_exceptionInfo_0_eSubCode <= stage1Out_thrown_payload_exceptionInfo_0_eSubCode;
      stage1Out_thrown_rData_exceptionInfo_1_exception <= stage1Out_thrown_payload_exceptionInfo_1_exception;
      stage1Out_thrown_rData_exceptionInfo_1_eCode <= stage1Out_thrown_payload_exceptionInfo_1_eCode;
      stage1Out_thrown_rData_exceptionInfo_1_eSubCode <= stage1Out_thrown_payload_exceptionInfo_1_eSubCode;
      stage1Out_thrown_rData_pc_0 <= stage1Out_thrown_payload_pc_0;
      stage1Out_thrown_rData_pc_1 <= stage1Out_thrown_payload_pc_1;
      stage1Out_thrown_rData_valid <= stage1Out_thrown_payload_valid;
      stage1Out_thrown_rData_tlb_hit <= stage1Out_thrown_payload_tlb_hit;
      stage1Out_thrown_rData_tlb_pageInfo_ppn <= stage1Out_thrown_payload_tlb_pageInfo_ppn;
      stage1Out_thrown_rData_tlb_pageInfo_plv <= stage1Out_thrown_payload_tlb_pageInfo_plv;
      stage1Out_thrown_rData_tlb_pageInfo_mat <= stage1Out_thrown_payload_tlb_pageInfo_mat;
      stage1Out_thrown_rData_tlb_pageInfo_d <= stage1Out_thrown_payload_tlb_pageInfo_d;
      stage1Out_thrown_rData_tlb_pageInfo_v <= stage1Out_thrown_payload_tlb_pageInfo_v;
      stage1Out_thrown_rData_wayValid_0 <= stage1Out_thrown_payload_wayValid_0;
      stage1Out_thrown_rData_wayValid_1 <= stage1Out_thrown_payload_wayValid_1;
      stage1Out_thrown_rData_isStoreTag <= stage1Out_thrown_payload_isStoreTag;
      stage1Out_thrown_rData_isIndexInvalidate <= stage1Out_thrown_payload_isIndexInvalidate;
      stage1Out_thrown_rData_isHitInvalidate <= stage1Out_thrown_payload_isHitInvalidate;
    end
    if(stage1Out_fire) begin
      fetchMask_0 <= 1'b0;
      fetchMask_1 <= 1'b0;
    end else begin
      fetchMask_0 <= (fetchMask_0 || bufWriteMask[0]);
    end
    if(stage1Out_fire) begin
      fetchMask_0 <= 1'b0;
      fetchMask_1 <= 1'b0;
    end else begin
      fetchMask_1 <= (fetchMask_1 || bufWriteMask[1]);
    end
    if(stage1Out_fire) begin
      wayOfReplace_0 <= 4'b0000;
    end
    if(stage1Out_fire) begin
      wayOfReplace_1 <= 4'b0000;
    end
    if(when_Cache_l255) begin
      missBuffer_0 <= io_axi_rdata;
    end
    if(when_Cache_l255_1) begin
      missBuffer_1 <= io_axi_rdata;
    end
    case(fsm_stateReg)
      fsm_enumDef_1_idle : begin
      end
      fsm_enumDef_1_req : begin
      end
      fsm_enumDef_1_read : begin
        if(when_Cache_l198) begin
          if(when_Cache_l200) begin
            transferBlockOffset <= (transferBlockOffset + 6'h04);
          end
          if(when_Cache_l200_1) begin
            transferBlockOffset <= (transferBlockOffset + 6'h04);
          end
          if(when_Cache_l200_2) begin
            transferBlockOffset <= (transferBlockOffset + 6'h04);
          end
          if(when_Cache_l200_3) begin
            transferBlockOffset <= (transferBlockOffset + 6'h04);
          end
        end
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l253) begin
      transferIndexOffset <= missAddr[11 : 6];
      transferBlockOffset <= missAddr[5 : 0];
      transferTag <= stage2In_payload_tlb_pageInfo_ppn;
      transferUncached <= (stage2In_payload_tlb_pageInfo_mat == 2'b00);
      replacingWay <= (_zz_missAddr ? wayToReplace_0 : wayToReplace_1);
    end
    if(when_StateMachine_l253_1) begin
      if(when_Cache_l180) begin
        if(when_Cache_l188) begin
          wayOfReplace_0 <= replacingWay;
        end
        if(when_Cache_l188_1) begin
          wayOfReplace_1 <= replacingWay;
        end
      end
    end
  end


endmodule

module NextLinePredictor (
  input  wire          io_pc_0_valid,
  input  wire [31:0]   io_pc_0_payload,
  input  wire          io_pc_1_valid,
  input  wire [31:0]   io_pc_1_payload,
  output wire          io_npc_0_valid,
  output wire [31:0]   io_npc_0_payload,
  output wire          io_npc_1_valid,
  output wire [31:0]   io_npc_1_payload,
  output wire [31:0]   io_branchInfo_0_predictPC,
  output wire          io_branchInfo_0_predictResult,
  output wire [31:0]   io_branchInfo_1_predictPC,
  output wire          io_branchInfo_1_predictResult,
  input  wire          io_updateInfo_0_valid,
  input  wire [31:0]   io_updateInfo_0_payload_pc,
  input  wire          io_updateInfo_0_payload_isJumpInst,
  input  wire          io_updateInfo_0_payload_taken,
  input  wire          io_updateInfo_0_payload_predictFail,
  input  wire [31:0]   io_updateInfo_0_payload_target,
  input  wire          io_updateInfo_1_valid,
  input  wire [31:0]   io_updateInfo_1_payload_pc,
  input  wire          io_updateInfo_1_payload_isJumpInst,
  input  wire          io_updateInfo_1_payload_taken,
  input  wire          io_updateInfo_1_payload_predictFail,
  input  wire [31:0]   io_updateInfo_1_payload_target
);

  wire       [1:0]    _zz__zz_lastPCIdx_2;
  reg        [31:0]   _zz_nextBase;
  reg        [1:0]    fetchMask;
  wire       [31:0]   nextBase;
  wire       [0:0]    lastPCIdx;
  wire       [1:0]    _zz_lastPCIdx;
  reg        [1:0]    _zz_lastPCIdx_1;
  wire       [1:0]    _zz_lastPCIdx_2;
  reg        [1:0]    _zz_lastPCIdx_3;
  wire                _zz_lastPCIdx_4;

  assign _zz__zz_lastPCIdx_2 = (_zz_lastPCIdx_1 - 2'b01);
  always @(*) begin
    case(lastPCIdx)
      1'b0 : _zz_nextBase = io_pc_0_payload;
      default : _zz_nextBase = io_pc_1_payload;
    endcase
  end

  assign _zz_lastPCIdx = fetchMask;
  always @(*) begin
    _zz_lastPCIdx_1[0] = _zz_lastPCIdx[1];
    _zz_lastPCIdx_1[1] = _zz_lastPCIdx[0];
  end

  assign _zz_lastPCIdx_2 = (_zz_lastPCIdx_1 & (~ _zz__zz_lastPCIdx_2));
  always @(*) begin
    _zz_lastPCIdx_3[0] = _zz_lastPCIdx_2[1];
    _zz_lastPCIdx_3[1] = _zz_lastPCIdx_2[0];
  end

  assign _zz_lastPCIdx_4 = _zz_lastPCIdx_3[1];
  assign lastPCIdx = _zz_lastPCIdx_4;
  assign nextBase = (_zz_nextBase + 32'h00000004);
  always @(*) begin
    fetchMask[0] = io_pc_0_valid;
    fetchMask[1] = io_pc_1_valid;
  end

  assign io_npc_0_valid = 1'b1;
  assign io_npc_0_payload = (nextBase + 32'h00000000);
  assign io_branchInfo_0_predictPC = 32'h00000000;
  assign io_branchInfo_0_predictResult = 1'b0;
  assign io_npc_1_valid = 1'b1;
  assign io_npc_1_payload = (nextBase + 32'h00000004);
  assign io_branchInfo_1_predictPC = 32'h00000000;
  assign io_branchInfo_1_predictResult = 1'b0;

endmodule

module PC (
  output wire          io_iCacheFeed_0_valid,
  input  wire          io_iCacheFeed_0_ready,
  output wire [31:0]   io_iCacheFeed_0_payload_address,
  output wire [3:0]    io_iCacheFeed_0_payload_size,
  output wire [31:0]   io_iCacheFeed_0_payload_branchInfo_predictPC,
  output wire          io_iCacheFeed_0_payload_branchInfo_predictResult,
  output wire          io_iCacheFeed_1_valid,
  input  wire          io_iCacheFeed_1_ready,
  output wire [31:0]   io_iCacheFeed_1_payload_address,
  output wire [3:0]    io_iCacheFeed_1_payload_size,
  output wire [31:0]   io_iCacheFeed_1_payload_branchInfo_predictPC,
  output wire          io_iCacheFeed_1_payload_branchInfo_predictResult,
  output wire          io_pc_0_valid,
  output wire [31:0]   io_pc_0_payload,
  output wire          io_pc_1_valid,
  output wire [31:0]   io_pc_1_payload,
  input  wire          io_npc_0_valid,
  input  wire [31:0]   io_npc_0_payload,
  input  wire          io_npc_1_valid,
  input  wire [31:0]   io_npc_1_payload,
  input  wire [31:0]   io_branchInfo_0_predictPC,
  input  wire          io_branchInfo_0_predictResult,
  input  wire [31:0]   io_branchInfo_1_predictPC,
  input  wire          io_branchInfo_1_predictResult,
  input  wire          io_flush,
  input  wire [31:0]   io_redirectPC,
  input  wire          aclk,
  input  wire          aresetn
);
  localparam LSUSizeOp_byte_1 = 4'd1;
  localparam LSUSizeOp_halfword = 4'd3;
  localparam LSUSizeOp_word = 4'd15;

  wire       [31:0]   _zz_pc_0_2;
  reg        [31:0]   _zz_pc_0_3;
  wire       [1:0]    _zz_pc_0_4;
  reg        [1:0]    _zz_pc_0_5;
  wire       [1:0]    _zz_pc_0_6;
  reg        [1:0]    _zz__zz_branchInfo_0_predictPC;
  wire       [1:0]    _zz__zz_branchInfo_0_predictPC_1;
  reg        [31:0]   _zz_branchInfo_0_predictPC_1;
  reg                 _zz_branchInfo_0_predictResult;
  reg                 _zz_valid_0;
  wire       [1:0]    _zz_valid_0_1;
  reg        [1:0]    _zz_valid_0_2;
  wire       [1:0]    _zz_valid_0_3;
  wire       [3:0]    _zz_nextPCListMid_1_0;
  wire       [3:0]    _zz__zz_nextBranchInfoListMid_1_0_predictPC;
  wire       [3:0]    _zz_nextValidListMid_1_0;
  wire       [3:0]    _zz_nextPCListMid_1_2;
  wire       [3:0]    _zz__zz_nextBranchInfoListMid_1_2_predictPC;
  wire       [3:0]    _zz_nextValidListMid_1_2;
  wire       [3:0]    _zz_nextPCListMid_1_1;
  wire       [3:0]    _zz__zz_nextBranchInfoListMid_1_1_predictPC;
  wire       [3:0]    _zz_nextValidListMid_1_1;
  wire       [3:0]    _zz_nextPCListMid_1_3;
  wire       [3:0]    _zz__zz_nextBranchInfoListMid_1_3_predictPC;
  wire       [3:0]    _zz_nextValidListMid_1_3;
  wire       [31:0]   _zz_pc_1;
  reg        [31:0]   _zz_pc_1_1;
  wire       [1:0]    _zz_pc_1_2;
  reg        [1:0]    _zz_pc_1_3;
  wire       [1:0]    _zz_pc_1_4;
  reg        [1:0]    _zz__zz_branchInfo_1_predictPC;
  wire       [1:0]    _zz__zz_branchInfo_1_predictPC_1;
  reg        [31:0]   _zz_branchInfo_1_predictPC_1;
  reg                 _zz_branchInfo_1_predictResult;
  reg                 _zz_valid_1;
  wire       [1:0]    _zz_valid_1_1;
  reg        [1:0]    _zz_valid_1_2;
  wire       [1:0]    _zz_valid_1_3;
  reg        [1:0]    acceptMask;
  reg        [31:0]   pc_0;
  reg        [31:0]   pc_1;
  reg        [31:0]   branchInfo_0_predictPC;
  reg                 branchInfo_0_predictResult;
  reg        [31:0]   branchInfo_1_predictPC;
  reg                 branchInfo_1_predictResult;
  reg                 valid_0;
  reg                 valid_1;
  wire       [31:0]   nextPCListMid_0_0;
  wire       [31:0]   nextPCListMid_0_1;
  wire       [31:0]   nextPCListMid_0_2;
  wire       [31:0]   nextPCListMid_0_3;
  wire       [31:0]   nextPCListMid_1_0;
  wire       [31:0]   nextPCListMid_1_1;
  wire       [31:0]   nextPCListMid_1_2;
  wire       [31:0]   nextPCListMid_1_3;
  wire       [31:0]   nextBranchInfoListMid_0_0_predictPC;
  wire                nextBranchInfoListMid_0_0_predictResult;
  wire       [31:0]   nextBranchInfoListMid_0_1_predictPC;
  wire                nextBranchInfoListMid_0_1_predictResult;
  wire       [31:0]   nextBranchInfoListMid_0_2_predictPC;
  wire                nextBranchInfoListMid_0_2_predictResult;
  wire       [31:0]   nextBranchInfoListMid_0_3_predictPC;
  wire                nextBranchInfoListMid_0_3_predictResult;
  wire       [31:0]   nextBranchInfoListMid_1_0_predictPC;
  wire                nextBranchInfoListMid_1_0_predictResult;
  wire       [31:0]   nextBranchInfoListMid_1_1_predictPC;
  wire                nextBranchInfoListMid_1_1_predictResult;
  wire       [31:0]   nextBranchInfoListMid_1_2_predictPC;
  wire                nextBranchInfoListMid_1_2_predictResult;
  wire       [31:0]   nextBranchInfoListMid_1_3_predictPC;
  wire                nextBranchInfoListMid_1_3_predictResult;
  wire                nextValidListMid_0_0;
  wire                nextValidListMid_0_1;
  wire                nextValidListMid_0_2;
  wire                nextValidListMid_0_3;
  wire                nextValidListMid_1_0;
  wire                nextValidListMid_1_1;
  wire                nextValidListMid_1_2;
  wire                nextValidListMid_1_3;
  wire       [31:0]   nextPCList_0;
  wire       [31:0]   nextPCList_1;
  wire       [31:0]   nextPCList_2;
  wire       [31:0]   nextPCList_3;
  wire       [31:0]   nextBranchInfoList_0_predictPC;
  wire                nextBranchInfoList_0_predictResult;
  wire       [31:0]   nextBranchInfoList_1_predictPC;
  wire                nextBranchInfoList_1_predictResult;
  wire       [31:0]   nextBranchInfoList_2_predictPC;
  wire                nextBranchInfoList_2_predictResult;
  wire       [31:0]   nextBranchInfoList_3_predictPC;
  wire                nextBranchInfoList_3_predictResult;
  wire                nextValidList_0;
  wire                nextValidList_1;
  wire                nextValidList_2;
  wire                nextValidList_3;
  wire                _zz_pc_0;
  wire                _zz_pc_0_1;
  wire       [1:0]    _zz_branchInfo_0_predictPC;
  wire                _zz_nextBranchInfoListMid_1_0_predictPC;
  wire                _zz_nextBranchInfoListMid_1_2_predictPC;
  wire                _zz_nextBranchInfoListMid_1_1_predictPC;
  wire                _zz_nextBranchInfoListMid_1_3_predictPC;
  wire       [1:0]    _zz_branchInfo_1_predictPC;
  `ifndef SYNTHESIS
  reg [63:0] io_iCacheFeed_0_payload_size_string;
  reg [63:0] io_iCacheFeed_1_payload_size_string;
  `endif


  assign _zz_pc_0_2 = (io_redirectPC + 32'h00000000);
  assign _zz_pc_0_4 = (2'b00 + _zz_pc_0_5);
  assign _zz_valid_0_1 = (2'b00 + _zz_valid_0_2);
  assign _zz_nextPCListMid_1_0 = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz__zz_nextBranchInfoListMid_1_0_predictPC = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz_nextValidListMid_1_0 = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz_nextPCListMid_1_2 = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz__zz_nextBranchInfoListMid_1_2_predictPC = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz_nextValidListMid_1_2 = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz_nextPCListMid_1_1 = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz__zz_nextBranchInfoListMid_1_1_predictPC = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz_nextValidListMid_1_1 = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz_nextPCListMid_1_3 = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz__zz_nextBranchInfoListMid_1_3_predictPC = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz_nextValidListMid_1_3 = {nextValidListMid_0_3,{nextValidListMid_0_2,{nextValidListMid_0_1,nextValidListMid_0_0}}};
  assign _zz_pc_1 = (io_redirectPC + 32'h00000004);
  assign _zz_pc_1_2 = (2'b01 + _zz_pc_1_3);
  assign _zz_valid_1_1 = (2'b01 + _zz_valid_1_2);
  assign _zz_pc_0_6 = {_zz_pc_0_1,_zz_pc_0};
  assign _zz__zz_branchInfo_0_predictPC_1 = {_zz_pc_0_1,_zz_pc_0};
  assign _zz_valid_0_3 = {_zz_pc_0_1,_zz_pc_0};
  assign _zz_pc_1_4 = {_zz_pc_0_1,_zz_pc_0};
  assign _zz__zz_branchInfo_1_predictPC_1 = {_zz_pc_0_1,_zz_pc_0};
  assign _zz_valid_1_3 = {_zz_pc_0_1,_zz_pc_0};
  always @(*) begin
    case(_zz_pc_0_4)
      2'b00 : _zz_pc_0_3 = nextPCListMid_1_0;
      2'b01 : _zz_pc_0_3 = nextPCListMid_1_1;
      2'b10 : _zz_pc_0_3 = nextPCListMid_1_2;
      default : _zz_pc_0_3 = nextPCListMid_1_3;
    endcase
  end

  always @(*) begin
    case(_zz_pc_0_6)
      2'b00 : _zz_pc_0_5 = 2'b00;
      2'b01 : _zz_pc_0_5 = 2'b01;
      2'b10 : _zz_pc_0_5 = 2'b01;
      default : _zz_pc_0_5 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz__zz_branchInfo_0_predictPC_1)
      2'b00 : _zz__zz_branchInfo_0_predictPC = 2'b00;
      2'b01 : _zz__zz_branchInfo_0_predictPC = 2'b01;
      2'b10 : _zz__zz_branchInfo_0_predictPC = 2'b01;
      default : _zz__zz_branchInfo_0_predictPC = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_branchInfo_0_predictPC)
      2'b00 : begin
        _zz_branchInfo_0_predictPC_1 = nextBranchInfoListMid_1_0_predictPC;
        _zz_branchInfo_0_predictResult = nextBranchInfoListMid_1_0_predictResult;
      end
      2'b01 : begin
        _zz_branchInfo_0_predictPC_1 = nextBranchInfoListMid_1_1_predictPC;
        _zz_branchInfo_0_predictResult = nextBranchInfoListMid_1_1_predictResult;
      end
      2'b10 : begin
        _zz_branchInfo_0_predictPC_1 = nextBranchInfoListMid_1_2_predictPC;
        _zz_branchInfo_0_predictResult = nextBranchInfoListMid_1_2_predictResult;
      end
      default : begin
        _zz_branchInfo_0_predictPC_1 = nextBranchInfoListMid_1_3_predictPC;
        _zz_branchInfo_0_predictResult = nextBranchInfoListMid_1_3_predictResult;
      end
    endcase
  end

  always @(*) begin
    case(_zz_valid_0_1)
      2'b00 : _zz_valid_0 = nextValidListMid_1_0;
      2'b01 : _zz_valid_0 = nextValidListMid_1_1;
      2'b10 : _zz_valid_0 = nextValidListMid_1_2;
      default : _zz_valid_0 = nextValidListMid_1_3;
    endcase
  end

  always @(*) begin
    case(_zz_valid_0_3)
      2'b00 : _zz_valid_0_2 = 2'b00;
      2'b01 : _zz_valid_0_2 = 2'b01;
      2'b10 : _zz_valid_0_2 = 2'b01;
      default : _zz_valid_0_2 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_pc_1_2)
      2'b00 : _zz_pc_1_1 = nextPCListMid_1_0;
      2'b01 : _zz_pc_1_1 = nextPCListMid_1_1;
      2'b10 : _zz_pc_1_1 = nextPCListMid_1_2;
      default : _zz_pc_1_1 = nextPCListMid_1_3;
    endcase
  end

  always @(*) begin
    case(_zz_pc_1_4)
      2'b00 : _zz_pc_1_3 = 2'b00;
      2'b01 : _zz_pc_1_3 = 2'b01;
      2'b10 : _zz_pc_1_3 = 2'b01;
      default : _zz_pc_1_3 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz__zz_branchInfo_1_predictPC_1)
      2'b00 : _zz__zz_branchInfo_1_predictPC = 2'b00;
      2'b01 : _zz__zz_branchInfo_1_predictPC = 2'b01;
      2'b10 : _zz__zz_branchInfo_1_predictPC = 2'b01;
      default : _zz__zz_branchInfo_1_predictPC = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_branchInfo_1_predictPC)
      2'b00 : begin
        _zz_branchInfo_1_predictPC_1 = nextBranchInfoListMid_1_0_predictPC;
        _zz_branchInfo_1_predictResult = nextBranchInfoListMid_1_0_predictResult;
      end
      2'b01 : begin
        _zz_branchInfo_1_predictPC_1 = nextBranchInfoListMid_1_1_predictPC;
        _zz_branchInfo_1_predictResult = nextBranchInfoListMid_1_1_predictResult;
      end
      2'b10 : begin
        _zz_branchInfo_1_predictPC_1 = nextBranchInfoListMid_1_2_predictPC;
        _zz_branchInfo_1_predictResult = nextBranchInfoListMid_1_2_predictResult;
      end
      default : begin
        _zz_branchInfo_1_predictPC_1 = nextBranchInfoListMid_1_3_predictPC;
        _zz_branchInfo_1_predictResult = nextBranchInfoListMid_1_3_predictResult;
      end
    endcase
  end

  always @(*) begin
    case(_zz_valid_1_1)
      2'b00 : _zz_valid_1 = nextValidListMid_1_0;
      2'b01 : _zz_valid_1 = nextValidListMid_1_1;
      2'b10 : _zz_valid_1 = nextValidListMid_1_2;
      default : _zz_valid_1 = nextValidListMid_1_3;
    endcase
  end

  always @(*) begin
    case(_zz_valid_1_3)
      2'b00 : _zz_valid_1_2 = 2'b00;
      2'b01 : _zz_valid_1_2 = 2'b01;
      2'b10 : _zz_valid_1_2 = 2'b01;
      default : _zz_valid_1_2 = 2'b10;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_iCacheFeed_0_payload_size)
      LSUSizeOp_byte_1 : io_iCacheFeed_0_payload_size_string = "byte_1  ";
      LSUSizeOp_halfword : io_iCacheFeed_0_payload_size_string = "halfword";
      LSUSizeOp_word : io_iCacheFeed_0_payload_size_string = "word    ";
      default : io_iCacheFeed_0_payload_size_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_iCacheFeed_1_payload_size)
      LSUSizeOp_byte_1 : io_iCacheFeed_1_payload_size_string = "byte_1  ";
      LSUSizeOp_halfword : io_iCacheFeed_1_payload_size_string = "halfword";
      LSUSizeOp_word : io_iCacheFeed_1_payload_size_string = "word    ";
      default : io_iCacheFeed_1_payload_size_string = "????????";
    endcase
  end
  `endif

  always @(*) begin
    acceptMask[0] = (io_iCacheFeed_0_ready && valid_0);
    acceptMask[1] = (io_iCacheFeed_1_ready && valid_1);
  end

  assign nextPCListMid_0_0 = pc_0;
  assign nextBranchInfoListMid_0_0_predictPC = branchInfo_0_predictPC;
  assign nextBranchInfoListMid_0_0_predictResult = branchInfo_0_predictResult;
  assign nextValidListMid_0_0 = valid_0;
  assign nextPCListMid_0_2 = io_npc_0_payload;
  assign nextValidListMid_0_2 = io_npc_0_valid;
  assign nextBranchInfoListMid_0_2_predictPC = io_branchInfo_0_predictPC;
  assign nextBranchInfoListMid_0_2_predictResult = io_branchInfo_0_predictResult;
  assign nextPCListMid_0_1 = pc_1;
  assign nextBranchInfoListMid_0_1_predictPC = branchInfo_1_predictPC;
  assign nextBranchInfoListMid_0_1_predictResult = branchInfo_1_predictResult;
  assign nextValidListMid_0_1 = valid_1;
  assign nextPCListMid_0_3 = io_npc_1_payload;
  assign nextValidListMid_0_3 = io_npc_1_valid;
  assign nextBranchInfoListMid_0_3_predictPC = io_branchInfo_1_predictPC;
  assign nextBranchInfoListMid_0_3_predictResult = io_branchInfo_1_predictResult;
  assign _zz_pc_0 = acceptMask[0];
  assign _zz_pc_0_1 = acceptMask[1];
  assign _zz_branchInfo_0_predictPC = (2'b00 + _zz__zz_branchInfo_0_predictPC);
  assign nextPCListMid_1_0 = ((&_zz_nextPCListMid_1_0[0 : 0]) ? nextPCListMid_0_0 : nextPCListMid_0_1);
  assign _zz_nextBranchInfoListMid_1_0_predictPC = (&_zz__zz_nextBranchInfoListMid_1_0_predictPC[0 : 0]);
  assign nextBranchInfoListMid_1_0_predictPC = (_zz_nextBranchInfoListMid_1_0_predictPC ? nextBranchInfoListMid_0_0_predictPC : nextBranchInfoListMid_0_1_predictPC);
  assign nextBranchInfoListMid_1_0_predictResult = (_zz_nextBranchInfoListMid_1_0_predictPC ? nextBranchInfoListMid_0_0_predictResult : nextBranchInfoListMid_0_1_predictResult);
  assign nextValidListMid_1_0 = ((&_zz_nextValidListMid_1_0[0 : 0]) ? nextValidListMid_0_0 : nextValidListMid_0_1);
  assign nextPCListMid_1_2 = ((&_zz_nextPCListMid_1_2[2 : 0]) ? nextPCListMid_0_2 : nextPCListMid_0_3);
  assign _zz_nextBranchInfoListMid_1_2_predictPC = (&_zz__zz_nextBranchInfoListMid_1_2_predictPC[2 : 0]);
  assign nextBranchInfoListMid_1_2_predictPC = (_zz_nextBranchInfoListMid_1_2_predictPC ? nextBranchInfoListMid_0_2_predictPC : nextBranchInfoListMid_0_3_predictPC);
  assign nextBranchInfoListMid_1_2_predictResult = (_zz_nextBranchInfoListMid_1_2_predictPC ? nextBranchInfoListMid_0_2_predictResult : nextBranchInfoListMid_0_3_predictResult);
  assign nextValidListMid_1_2 = ((&_zz_nextValidListMid_1_2[2 : 0]) ? nextValidListMid_0_2 : nextValidListMid_0_3);
  assign nextPCListMid_1_1 = ((&_zz_nextPCListMid_1_1[1 : 0]) ? nextPCListMid_0_1 : nextPCListMid_0_2);
  assign _zz_nextBranchInfoListMid_1_1_predictPC = (&_zz__zz_nextBranchInfoListMid_1_1_predictPC[1 : 0]);
  assign nextBranchInfoListMid_1_1_predictPC = (_zz_nextBranchInfoListMid_1_1_predictPC ? nextBranchInfoListMid_0_1_predictPC : nextBranchInfoListMid_0_2_predictPC);
  assign nextBranchInfoListMid_1_1_predictResult = (_zz_nextBranchInfoListMid_1_1_predictPC ? nextBranchInfoListMid_0_1_predictResult : nextBranchInfoListMid_0_2_predictResult);
  assign nextValidListMid_1_1 = ((&_zz_nextValidListMid_1_1[1 : 0]) ? nextValidListMid_0_1 : nextValidListMid_0_2);
  assign nextPCListMid_1_3 = ((&_zz_nextPCListMid_1_3[3 : 0]) ? nextPCListMid_0_3 : 32'h00000000);
  assign _zz_nextBranchInfoListMid_1_3_predictPC = (&_zz__zz_nextBranchInfoListMid_1_3_predictPC[3 : 0]);
  assign nextBranchInfoListMid_1_3_predictPC = (_zz_nextBranchInfoListMid_1_3_predictPC ? nextBranchInfoListMid_0_3_predictPC : 32'h00000000);
  assign nextBranchInfoListMid_1_3_predictResult = (_zz_nextBranchInfoListMid_1_3_predictPC ? nextBranchInfoListMid_0_3_predictResult : 1'b0);
  assign nextValidListMid_1_3 = ((&_zz_nextValidListMid_1_3[3 : 0]) ? nextValidListMid_0_3 : 1'b0);
  assign _zz_branchInfo_1_predictPC = (2'b01 + _zz__zz_branchInfo_1_predictPC);
  assign io_iCacheFeed_0_valid = valid_0;
  assign io_iCacheFeed_0_payload_address = pc_0;
  assign io_iCacheFeed_0_payload_size = LSUSizeOp_word;
  assign io_iCacheFeed_0_payload_branchInfo_predictPC = branchInfo_0_predictPC;
  assign io_iCacheFeed_0_payload_branchInfo_predictResult = branchInfo_0_predictResult;
  assign io_pc_0_valid = valid_0;
  assign io_pc_0_payload = pc_0;
  assign io_iCacheFeed_1_valid = valid_1;
  assign io_iCacheFeed_1_payload_address = pc_1;
  assign io_iCacheFeed_1_payload_size = LSUSizeOp_word;
  assign io_iCacheFeed_1_payload_branchInfo_predictPC = branchInfo_1_predictPC;
  assign io_iCacheFeed_1_payload_branchInfo_predictResult = branchInfo_1_predictResult;
  assign io_pc_1_valid = valid_1;
  assign io_pc_1_payload = pc_1;
  always @(posedge aclk) begin
    if(!aresetn) begin
      pc_0 <= 32'h1c000000;
      branchInfo_0_predictPC <= 32'h00000000;
      branchInfo_0_predictResult <= 1'b0;
      valid_0 <= 1'b1;
      pc_1 <= 32'h1c000004;
      branchInfo_1_predictPC <= 32'h00000000;
      branchInfo_1_predictResult <= 1'b0;
      valid_1 <= 1'b1;
    end else begin
      pc_0 <= (io_flush ? _zz_pc_0_2 : _zz_pc_0_3);
      branchInfo_0_predictPC <= (io_flush ? 32'h00000000 : _zz_branchInfo_0_predictPC_1);
      branchInfo_0_predictResult <= (io_flush ? 1'b0 : _zz_branchInfo_0_predictResult);
      valid_0 <= (io_flush ? 1'b1 : _zz_valid_0);
      pc_1 <= (io_flush ? _zz_pc_1 : _zz_pc_1_1);
      branchInfo_1_predictPC <= (io_flush ? 32'h00000000 : _zz_branchInfo_1_predictPC_1);
      branchInfo_1_predictResult <= (io_flush ? 1'b0 : _zz_branchInfo_1_predictResult);
      valid_1 <= (io_flush ? 1'b1 : _zz_valid_1);
    end
  end


endmodule

module FreeList (
  input  wire [1:0]    io_dispatch_disPatchNum,
  output reg  [1:0]    io_dispatch_availMask,
  output wire [5:0]    io_dispatch_prfIdx_0,
  output wire [5:0]    io_dispatch_prfIdx_1,
  input  wire [5:0]    io_retire_prfIdx_0,
  input  wire [5:0]    io_retire_prfIdx_1,
  input  wire [1:0]    io_retire_writeNum,
  input  wire          io_retire_delayedFlush,
  input  wire          aclk,
  input  wire          aresetn
);

  wire       [0:0]    _zz_retirePtr;
  reg        [5:0]    _zz_io_dispatch_prfIdx_0;
  wire       [5:0]    _zz_allocPtr_0;
  reg        [5:0]    _zz_io_dispatch_prfIdx_1;
  wire       [5:0]    _zz_allocPtr_1;
  wire       [0:0]    _zz_retireEnableMask;
  wire       [5:0]    _zz_freePtr_0;
  wire       [5:0]    _zz_freePtr_1;
  wire       [5:0]    _zz_retirePtr_1;
  reg        [5:0]    freeList_0;
  reg        [5:0]    freeList_1;
  reg        [5:0]    freeList_2;
  reg        [5:0]    freeList_3;
  reg        [5:0]    freeList_4;
  reg        [5:0]    freeList_5;
  reg        [5:0]    freeList_6;
  reg        [5:0]    freeList_7;
  reg        [5:0]    freeList_8;
  reg        [5:0]    freeList_9;
  reg        [5:0]    freeList_10;
  reg        [5:0]    freeList_11;
  reg        [5:0]    freeList_12;
  reg        [5:0]    freeList_13;
  reg        [5:0]    freeList_14;
  reg        [5:0]    freeList_15;
  reg        [5:0]    freeList_16;
  reg        [5:0]    freeList_17;
  reg        [5:0]    freeList_18;
  reg        [5:0]    freeList_19;
  reg        [5:0]    freeList_20;
  reg        [5:0]    freeList_21;
  reg        [5:0]    freeList_22;
  reg        [5:0]    freeList_23;
  reg        [5:0]    freeList_24;
  reg        [5:0]    freeList_25;
  reg        [5:0]    freeList_26;
  reg        [5:0]    freeList_27;
  reg        [5:0]    freeList_28;
  reg        [5:0]    freeList_29;
  reg        [5:0]    freeList_30;
  reg        [5:0]    freeList_31;
  reg        [5:0]    freeList_32;
  reg        [5:0]    freeList_33;
  reg        [5:0]    freeList_34;
  reg        [5:0]    freeList_35;
  reg        [5:0]    freeList_36;
  reg        [5:0]    freeList_37;
  reg        [5:0]    freeList_38;
  reg        [5:0]    freeList_39;
  reg        [5:0]    freeList_40;
  reg        [5:0]    freeList_41;
  reg        [5:0]    freeList_42;
  reg        [5:0]    freeList_43;
  reg        [5:0]    freeList_44;
  reg        [5:0]    freeList_45;
  reg        [5:0]    freeList_46;
  reg        [5:0]    freeList_47;
  reg        [5:0]    freeList_48;
  reg        [5:0]    freeList_49;
  reg        [5:0]    freeList_50;
  reg        [5:0]    freeList_51;
  reg        [5:0]    freeList_52;
  reg        [5:0]    freeList_53;
  reg        [5:0]    freeList_54;
  reg        [5:0]    freeList_55;
  reg        [5:0]    freeList_56;
  reg        [5:0]    freeList_57;
  reg        [5:0]    freeList_58;
  reg        [5:0]    freeList_59;
  reg        [5:0]    freeList_60;
  reg        [5:0]    freeList_61;
  reg        [5:0]    freeList_62;
  reg        [5:0]    freeList_63;
  reg        [5:0]    freePtr_0;
  reg        [5:0]    freePtr_1;
  reg        [5:0]    allocPtr_0;
  reg        [5:0]    allocPtr_1;
  reg        [5:0]    retirePtr;
  reg        [1:0]    availMask;
  reg        [1:0]    retireEnableMask;
  wire                when_RAT_l101;
  wire       [63:0]   _zz_1;
  wire                when_RAT_l101_1;
  wire       [63:0]   _zz_2;

  assign _zz_retirePtr = 1'b1;
  assign _zz_allocPtr_0 = {4'd0, io_dispatch_disPatchNum};
  assign _zz_allocPtr_1 = {4'd0, io_dispatch_disPatchNum};
  assign _zz_retireEnableMask = 1'b1;
  assign _zz_freePtr_0 = {4'd0, io_retire_writeNum};
  assign _zz_freePtr_1 = {4'd0, io_retire_writeNum};
  assign _zz_retirePtr_1 = {4'd0, io_retire_writeNum};
  always @(*) begin
    case(allocPtr_0)
      6'b000000 : _zz_io_dispatch_prfIdx_0 = freeList_0;
      6'b000001 : _zz_io_dispatch_prfIdx_0 = freeList_1;
      6'b000010 : _zz_io_dispatch_prfIdx_0 = freeList_2;
      6'b000011 : _zz_io_dispatch_prfIdx_0 = freeList_3;
      6'b000100 : _zz_io_dispatch_prfIdx_0 = freeList_4;
      6'b000101 : _zz_io_dispatch_prfIdx_0 = freeList_5;
      6'b000110 : _zz_io_dispatch_prfIdx_0 = freeList_6;
      6'b000111 : _zz_io_dispatch_prfIdx_0 = freeList_7;
      6'b001000 : _zz_io_dispatch_prfIdx_0 = freeList_8;
      6'b001001 : _zz_io_dispatch_prfIdx_0 = freeList_9;
      6'b001010 : _zz_io_dispatch_prfIdx_0 = freeList_10;
      6'b001011 : _zz_io_dispatch_prfIdx_0 = freeList_11;
      6'b001100 : _zz_io_dispatch_prfIdx_0 = freeList_12;
      6'b001101 : _zz_io_dispatch_prfIdx_0 = freeList_13;
      6'b001110 : _zz_io_dispatch_prfIdx_0 = freeList_14;
      6'b001111 : _zz_io_dispatch_prfIdx_0 = freeList_15;
      6'b010000 : _zz_io_dispatch_prfIdx_0 = freeList_16;
      6'b010001 : _zz_io_dispatch_prfIdx_0 = freeList_17;
      6'b010010 : _zz_io_dispatch_prfIdx_0 = freeList_18;
      6'b010011 : _zz_io_dispatch_prfIdx_0 = freeList_19;
      6'b010100 : _zz_io_dispatch_prfIdx_0 = freeList_20;
      6'b010101 : _zz_io_dispatch_prfIdx_0 = freeList_21;
      6'b010110 : _zz_io_dispatch_prfIdx_0 = freeList_22;
      6'b010111 : _zz_io_dispatch_prfIdx_0 = freeList_23;
      6'b011000 : _zz_io_dispatch_prfIdx_0 = freeList_24;
      6'b011001 : _zz_io_dispatch_prfIdx_0 = freeList_25;
      6'b011010 : _zz_io_dispatch_prfIdx_0 = freeList_26;
      6'b011011 : _zz_io_dispatch_prfIdx_0 = freeList_27;
      6'b011100 : _zz_io_dispatch_prfIdx_0 = freeList_28;
      6'b011101 : _zz_io_dispatch_prfIdx_0 = freeList_29;
      6'b011110 : _zz_io_dispatch_prfIdx_0 = freeList_30;
      6'b011111 : _zz_io_dispatch_prfIdx_0 = freeList_31;
      6'b100000 : _zz_io_dispatch_prfIdx_0 = freeList_32;
      6'b100001 : _zz_io_dispatch_prfIdx_0 = freeList_33;
      6'b100010 : _zz_io_dispatch_prfIdx_0 = freeList_34;
      6'b100011 : _zz_io_dispatch_prfIdx_0 = freeList_35;
      6'b100100 : _zz_io_dispatch_prfIdx_0 = freeList_36;
      6'b100101 : _zz_io_dispatch_prfIdx_0 = freeList_37;
      6'b100110 : _zz_io_dispatch_prfIdx_0 = freeList_38;
      6'b100111 : _zz_io_dispatch_prfIdx_0 = freeList_39;
      6'b101000 : _zz_io_dispatch_prfIdx_0 = freeList_40;
      6'b101001 : _zz_io_dispatch_prfIdx_0 = freeList_41;
      6'b101010 : _zz_io_dispatch_prfIdx_0 = freeList_42;
      6'b101011 : _zz_io_dispatch_prfIdx_0 = freeList_43;
      6'b101100 : _zz_io_dispatch_prfIdx_0 = freeList_44;
      6'b101101 : _zz_io_dispatch_prfIdx_0 = freeList_45;
      6'b101110 : _zz_io_dispatch_prfIdx_0 = freeList_46;
      6'b101111 : _zz_io_dispatch_prfIdx_0 = freeList_47;
      6'b110000 : _zz_io_dispatch_prfIdx_0 = freeList_48;
      6'b110001 : _zz_io_dispatch_prfIdx_0 = freeList_49;
      6'b110010 : _zz_io_dispatch_prfIdx_0 = freeList_50;
      6'b110011 : _zz_io_dispatch_prfIdx_0 = freeList_51;
      6'b110100 : _zz_io_dispatch_prfIdx_0 = freeList_52;
      6'b110101 : _zz_io_dispatch_prfIdx_0 = freeList_53;
      6'b110110 : _zz_io_dispatch_prfIdx_0 = freeList_54;
      6'b110111 : _zz_io_dispatch_prfIdx_0 = freeList_55;
      6'b111000 : _zz_io_dispatch_prfIdx_0 = freeList_56;
      6'b111001 : _zz_io_dispatch_prfIdx_0 = freeList_57;
      6'b111010 : _zz_io_dispatch_prfIdx_0 = freeList_58;
      6'b111011 : _zz_io_dispatch_prfIdx_0 = freeList_59;
      6'b111100 : _zz_io_dispatch_prfIdx_0 = freeList_60;
      6'b111101 : _zz_io_dispatch_prfIdx_0 = freeList_61;
      6'b111110 : _zz_io_dispatch_prfIdx_0 = freeList_62;
      default : _zz_io_dispatch_prfIdx_0 = freeList_63;
    endcase
  end

  always @(*) begin
    case(allocPtr_1)
      6'b000000 : _zz_io_dispatch_prfIdx_1 = freeList_0;
      6'b000001 : _zz_io_dispatch_prfIdx_1 = freeList_1;
      6'b000010 : _zz_io_dispatch_prfIdx_1 = freeList_2;
      6'b000011 : _zz_io_dispatch_prfIdx_1 = freeList_3;
      6'b000100 : _zz_io_dispatch_prfIdx_1 = freeList_4;
      6'b000101 : _zz_io_dispatch_prfIdx_1 = freeList_5;
      6'b000110 : _zz_io_dispatch_prfIdx_1 = freeList_6;
      6'b000111 : _zz_io_dispatch_prfIdx_1 = freeList_7;
      6'b001000 : _zz_io_dispatch_prfIdx_1 = freeList_8;
      6'b001001 : _zz_io_dispatch_prfIdx_1 = freeList_9;
      6'b001010 : _zz_io_dispatch_prfIdx_1 = freeList_10;
      6'b001011 : _zz_io_dispatch_prfIdx_1 = freeList_11;
      6'b001100 : _zz_io_dispatch_prfIdx_1 = freeList_12;
      6'b001101 : _zz_io_dispatch_prfIdx_1 = freeList_13;
      6'b001110 : _zz_io_dispatch_prfIdx_1 = freeList_14;
      6'b001111 : _zz_io_dispatch_prfIdx_1 = freeList_15;
      6'b010000 : _zz_io_dispatch_prfIdx_1 = freeList_16;
      6'b010001 : _zz_io_dispatch_prfIdx_1 = freeList_17;
      6'b010010 : _zz_io_dispatch_prfIdx_1 = freeList_18;
      6'b010011 : _zz_io_dispatch_prfIdx_1 = freeList_19;
      6'b010100 : _zz_io_dispatch_prfIdx_1 = freeList_20;
      6'b010101 : _zz_io_dispatch_prfIdx_1 = freeList_21;
      6'b010110 : _zz_io_dispatch_prfIdx_1 = freeList_22;
      6'b010111 : _zz_io_dispatch_prfIdx_1 = freeList_23;
      6'b011000 : _zz_io_dispatch_prfIdx_1 = freeList_24;
      6'b011001 : _zz_io_dispatch_prfIdx_1 = freeList_25;
      6'b011010 : _zz_io_dispatch_prfIdx_1 = freeList_26;
      6'b011011 : _zz_io_dispatch_prfIdx_1 = freeList_27;
      6'b011100 : _zz_io_dispatch_prfIdx_1 = freeList_28;
      6'b011101 : _zz_io_dispatch_prfIdx_1 = freeList_29;
      6'b011110 : _zz_io_dispatch_prfIdx_1 = freeList_30;
      6'b011111 : _zz_io_dispatch_prfIdx_1 = freeList_31;
      6'b100000 : _zz_io_dispatch_prfIdx_1 = freeList_32;
      6'b100001 : _zz_io_dispatch_prfIdx_1 = freeList_33;
      6'b100010 : _zz_io_dispatch_prfIdx_1 = freeList_34;
      6'b100011 : _zz_io_dispatch_prfIdx_1 = freeList_35;
      6'b100100 : _zz_io_dispatch_prfIdx_1 = freeList_36;
      6'b100101 : _zz_io_dispatch_prfIdx_1 = freeList_37;
      6'b100110 : _zz_io_dispatch_prfIdx_1 = freeList_38;
      6'b100111 : _zz_io_dispatch_prfIdx_1 = freeList_39;
      6'b101000 : _zz_io_dispatch_prfIdx_1 = freeList_40;
      6'b101001 : _zz_io_dispatch_prfIdx_1 = freeList_41;
      6'b101010 : _zz_io_dispatch_prfIdx_1 = freeList_42;
      6'b101011 : _zz_io_dispatch_prfIdx_1 = freeList_43;
      6'b101100 : _zz_io_dispatch_prfIdx_1 = freeList_44;
      6'b101101 : _zz_io_dispatch_prfIdx_1 = freeList_45;
      6'b101110 : _zz_io_dispatch_prfIdx_1 = freeList_46;
      6'b101111 : _zz_io_dispatch_prfIdx_1 = freeList_47;
      6'b110000 : _zz_io_dispatch_prfIdx_1 = freeList_48;
      6'b110001 : _zz_io_dispatch_prfIdx_1 = freeList_49;
      6'b110010 : _zz_io_dispatch_prfIdx_1 = freeList_50;
      6'b110011 : _zz_io_dispatch_prfIdx_1 = freeList_51;
      6'b110100 : _zz_io_dispatch_prfIdx_1 = freeList_52;
      6'b110101 : _zz_io_dispatch_prfIdx_1 = freeList_53;
      6'b110110 : _zz_io_dispatch_prfIdx_1 = freeList_54;
      6'b110111 : _zz_io_dispatch_prfIdx_1 = freeList_55;
      6'b111000 : _zz_io_dispatch_prfIdx_1 = freeList_56;
      6'b111001 : _zz_io_dispatch_prfIdx_1 = freeList_57;
      6'b111010 : _zz_io_dispatch_prfIdx_1 = freeList_58;
      6'b111011 : _zz_io_dispatch_prfIdx_1 = freeList_59;
      6'b111100 : _zz_io_dispatch_prfIdx_1 = freeList_60;
      6'b111101 : _zz_io_dispatch_prfIdx_1 = freeList_61;
      6'b111110 : _zz_io_dispatch_prfIdx_1 = freeList_62;
      default : _zz_io_dispatch_prfIdx_1 = freeList_63;
    endcase
  end

  always @(*) begin
    availMask[0] = (allocPtr_0 != freePtr_0);
    availMask[1] = (allocPtr_1 != freePtr_0);
  end

  always @(*) begin
    io_dispatch_availMask[0] = (&availMask[0 : 0]);
    io_dispatch_availMask[1] = (&availMask[1 : 0]);
  end

  assign io_dispatch_prfIdx_0 = _zz_io_dispatch_prfIdx_0;
  assign io_dispatch_prfIdx_1 = _zz_io_dispatch_prfIdx_1;
  always @(*) begin
    retireEnableMask = 2'bxx;
    case(io_retire_writeNum)
      2'b00 : begin
        retireEnableMask = 2'b00;
      end
      2'b01 : begin
        retireEnableMask = {1'd0, _zz_retireEnableMask};
      end
      2'b10 : begin
        retireEnableMask = 2'b11;
      end
      default : begin
      end
    endcase
  end

  assign when_RAT_l101 = retireEnableMask[0];
  assign _zz_1 = ({63'd0,1'b1} <<< freePtr_0);
  assign when_RAT_l101_1 = retireEnableMask[1];
  assign _zz_2 = ({63'd0,1'b1} <<< freePtr_1);
  always @(posedge aclk) begin
    if(!aresetn) begin
      freeList_0 <= 6'h00;
      freeList_1 <= 6'h01;
      freeList_2 <= 6'h02;
      freeList_3 <= 6'h03;
      freeList_4 <= 6'h04;
      freeList_5 <= 6'h05;
      freeList_6 <= 6'h06;
      freeList_7 <= 6'h07;
      freeList_8 <= 6'h08;
      freeList_9 <= 6'h09;
      freeList_10 <= 6'h0a;
      freeList_11 <= 6'h0b;
      freeList_12 <= 6'h0c;
      freeList_13 <= 6'h0d;
      freeList_14 <= 6'h0e;
      freeList_15 <= 6'h0f;
      freeList_16 <= 6'h10;
      freeList_17 <= 6'h11;
      freeList_18 <= 6'h12;
      freeList_19 <= 6'h13;
      freeList_20 <= 6'h14;
      freeList_21 <= 6'h15;
      freeList_22 <= 6'h16;
      freeList_23 <= 6'h17;
      freeList_24 <= 6'h18;
      freeList_25 <= 6'h19;
      freeList_26 <= 6'h1a;
      freeList_27 <= 6'h1b;
      freeList_28 <= 6'h1c;
      freeList_29 <= 6'h1d;
      freeList_30 <= 6'h1e;
      freeList_31 <= 6'h1f;
      freeList_32 <= 6'h20;
      freeList_33 <= 6'h21;
      freeList_34 <= 6'h22;
      freeList_35 <= 6'h23;
      freeList_36 <= 6'h24;
      freeList_37 <= 6'h25;
      freeList_38 <= 6'h26;
      freeList_39 <= 6'h27;
      freeList_40 <= 6'h28;
      freeList_41 <= 6'h29;
      freeList_42 <= 6'h2a;
      freeList_43 <= 6'h2b;
      freeList_44 <= 6'h2c;
      freeList_45 <= 6'h2d;
      freeList_46 <= 6'h2e;
      freeList_47 <= 6'h2f;
      freeList_48 <= 6'h30;
      freeList_49 <= 6'h31;
      freeList_50 <= 6'h32;
      freeList_51 <= 6'h33;
      freeList_52 <= 6'h34;
      freeList_53 <= 6'h35;
      freeList_54 <= 6'h36;
      freeList_55 <= 6'h37;
      freeList_56 <= 6'h38;
      freeList_57 <= 6'h39;
      freeList_58 <= 6'h3a;
      freeList_59 <= 6'h3b;
      freeList_60 <= 6'h3c;
      freeList_61 <= 6'h3d;
      freeList_62 <= 6'h3e;
      freeList_63 <= 6'h3f;
      freePtr_0 <= 6'h00;
      freePtr_1 <= 6'h01;
      allocPtr_0 <= 6'h01;
      allocPtr_1 <= 6'h02;
      retirePtr <= {5'd0, _zz_retirePtr};
    end else begin
      allocPtr_0 <= (allocPtr_0 + _zz_allocPtr_0);
      allocPtr_1 <= (allocPtr_1 + _zz_allocPtr_1);
      if(when_RAT_l101) begin
        if(_zz_1[0]) begin
          freeList_0 <= io_retire_prfIdx_0;
        end
        if(_zz_1[1]) begin
          freeList_1 <= io_retire_prfIdx_0;
        end
        if(_zz_1[2]) begin
          freeList_2 <= io_retire_prfIdx_0;
        end
        if(_zz_1[3]) begin
          freeList_3 <= io_retire_prfIdx_0;
        end
        if(_zz_1[4]) begin
          freeList_4 <= io_retire_prfIdx_0;
        end
        if(_zz_1[5]) begin
          freeList_5 <= io_retire_prfIdx_0;
        end
        if(_zz_1[6]) begin
          freeList_6 <= io_retire_prfIdx_0;
        end
        if(_zz_1[7]) begin
          freeList_7 <= io_retire_prfIdx_0;
        end
        if(_zz_1[8]) begin
          freeList_8 <= io_retire_prfIdx_0;
        end
        if(_zz_1[9]) begin
          freeList_9 <= io_retire_prfIdx_0;
        end
        if(_zz_1[10]) begin
          freeList_10 <= io_retire_prfIdx_0;
        end
        if(_zz_1[11]) begin
          freeList_11 <= io_retire_prfIdx_0;
        end
        if(_zz_1[12]) begin
          freeList_12 <= io_retire_prfIdx_0;
        end
        if(_zz_1[13]) begin
          freeList_13 <= io_retire_prfIdx_0;
        end
        if(_zz_1[14]) begin
          freeList_14 <= io_retire_prfIdx_0;
        end
        if(_zz_1[15]) begin
          freeList_15 <= io_retire_prfIdx_0;
        end
        if(_zz_1[16]) begin
          freeList_16 <= io_retire_prfIdx_0;
        end
        if(_zz_1[17]) begin
          freeList_17 <= io_retire_prfIdx_0;
        end
        if(_zz_1[18]) begin
          freeList_18 <= io_retire_prfIdx_0;
        end
        if(_zz_1[19]) begin
          freeList_19 <= io_retire_prfIdx_0;
        end
        if(_zz_1[20]) begin
          freeList_20 <= io_retire_prfIdx_0;
        end
        if(_zz_1[21]) begin
          freeList_21 <= io_retire_prfIdx_0;
        end
        if(_zz_1[22]) begin
          freeList_22 <= io_retire_prfIdx_0;
        end
        if(_zz_1[23]) begin
          freeList_23 <= io_retire_prfIdx_0;
        end
        if(_zz_1[24]) begin
          freeList_24 <= io_retire_prfIdx_0;
        end
        if(_zz_1[25]) begin
          freeList_25 <= io_retire_prfIdx_0;
        end
        if(_zz_1[26]) begin
          freeList_26 <= io_retire_prfIdx_0;
        end
        if(_zz_1[27]) begin
          freeList_27 <= io_retire_prfIdx_0;
        end
        if(_zz_1[28]) begin
          freeList_28 <= io_retire_prfIdx_0;
        end
        if(_zz_1[29]) begin
          freeList_29 <= io_retire_prfIdx_0;
        end
        if(_zz_1[30]) begin
          freeList_30 <= io_retire_prfIdx_0;
        end
        if(_zz_1[31]) begin
          freeList_31 <= io_retire_prfIdx_0;
        end
        if(_zz_1[32]) begin
          freeList_32 <= io_retire_prfIdx_0;
        end
        if(_zz_1[33]) begin
          freeList_33 <= io_retire_prfIdx_0;
        end
        if(_zz_1[34]) begin
          freeList_34 <= io_retire_prfIdx_0;
        end
        if(_zz_1[35]) begin
          freeList_35 <= io_retire_prfIdx_0;
        end
        if(_zz_1[36]) begin
          freeList_36 <= io_retire_prfIdx_0;
        end
        if(_zz_1[37]) begin
          freeList_37 <= io_retire_prfIdx_0;
        end
        if(_zz_1[38]) begin
          freeList_38 <= io_retire_prfIdx_0;
        end
        if(_zz_1[39]) begin
          freeList_39 <= io_retire_prfIdx_0;
        end
        if(_zz_1[40]) begin
          freeList_40 <= io_retire_prfIdx_0;
        end
        if(_zz_1[41]) begin
          freeList_41 <= io_retire_prfIdx_0;
        end
        if(_zz_1[42]) begin
          freeList_42 <= io_retire_prfIdx_0;
        end
        if(_zz_1[43]) begin
          freeList_43 <= io_retire_prfIdx_0;
        end
        if(_zz_1[44]) begin
          freeList_44 <= io_retire_prfIdx_0;
        end
        if(_zz_1[45]) begin
          freeList_45 <= io_retire_prfIdx_0;
        end
        if(_zz_1[46]) begin
          freeList_46 <= io_retire_prfIdx_0;
        end
        if(_zz_1[47]) begin
          freeList_47 <= io_retire_prfIdx_0;
        end
        if(_zz_1[48]) begin
          freeList_48 <= io_retire_prfIdx_0;
        end
        if(_zz_1[49]) begin
          freeList_49 <= io_retire_prfIdx_0;
        end
        if(_zz_1[50]) begin
          freeList_50 <= io_retire_prfIdx_0;
        end
        if(_zz_1[51]) begin
          freeList_51 <= io_retire_prfIdx_0;
        end
        if(_zz_1[52]) begin
          freeList_52 <= io_retire_prfIdx_0;
        end
        if(_zz_1[53]) begin
          freeList_53 <= io_retire_prfIdx_0;
        end
        if(_zz_1[54]) begin
          freeList_54 <= io_retire_prfIdx_0;
        end
        if(_zz_1[55]) begin
          freeList_55 <= io_retire_prfIdx_0;
        end
        if(_zz_1[56]) begin
          freeList_56 <= io_retire_prfIdx_0;
        end
        if(_zz_1[57]) begin
          freeList_57 <= io_retire_prfIdx_0;
        end
        if(_zz_1[58]) begin
          freeList_58 <= io_retire_prfIdx_0;
        end
        if(_zz_1[59]) begin
          freeList_59 <= io_retire_prfIdx_0;
        end
        if(_zz_1[60]) begin
          freeList_60 <= io_retire_prfIdx_0;
        end
        if(_zz_1[61]) begin
          freeList_61 <= io_retire_prfIdx_0;
        end
        if(_zz_1[62]) begin
          freeList_62 <= io_retire_prfIdx_0;
        end
        if(_zz_1[63]) begin
          freeList_63 <= io_retire_prfIdx_0;
        end
      end
      freePtr_0 <= (freePtr_0 + _zz_freePtr_0);
      if(when_RAT_l101_1) begin
        if(_zz_2[0]) begin
          freeList_0 <= io_retire_prfIdx_1;
        end
        if(_zz_2[1]) begin
          freeList_1 <= io_retire_prfIdx_1;
        end
        if(_zz_2[2]) begin
          freeList_2 <= io_retire_prfIdx_1;
        end
        if(_zz_2[3]) begin
          freeList_3 <= io_retire_prfIdx_1;
        end
        if(_zz_2[4]) begin
          freeList_4 <= io_retire_prfIdx_1;
        end
        if(_zz_2[5]) begin
          freeList_5 <= io_retire_prfIdx_1;
        end
        if(_zz_2[6]) begin
          freeList_6 <= io_retire_prfIdx_1;
        end
        if(_zz_2[7]) begin
          freeList_7 <= io_retire_prfIdx_1;
        end
        if(_zz_2[8]) begin
          freeList_8 <= io_retire_prfIdx_1;
        end
        if(_zz_2[9]) begin
          freeList_9 <= io_retire_prfIdx_1;
        end
        if(_zz_2[10]) begin
          freeList_10 <= io_retire_prfIdx_1;
        end
        if(_zz_2[11]) begin
          freeList_11 <= io_retire_prfIdx_1;
        end
        if(_zz_2[12]) begin
          freeList_12 <= io_retire_prfIdx_1;
        end
        if(_zz_2[13]) begin
          freeList_13 <= io_retire_prfIdx_1;
        end
        if(_zz_2[14]) begin
          freeList_14 <= io_retire_prfIdx_1;
        end
        if(_zz_2[15]) begin
          freeList_15 <= io_retire_prfIdx_1;
        end
        if(_zz_2[16]) begin
          freeList_16 <= io_retire_prfIdx_1;
        end
        if(_zz_2[17]) begin
          freeList_17 <= io_retire_prfIdx_1;
        end
        if(_zz_2[18]) begin
          freeList_18 <= io_retire_prfIdx_1;
        end
        if(_zz_2[19]) begin
          freeList_19 <= io_retire_prfIdx_1;
        end
        if(_zz_2[20]) begin
          freeList_20 <= io_retire_prfIdx_1;
        end
        if(_zz_2[21]) begin
          freeList_21 <= io_retire_prfIdx_1;
        end
        if(_zz_2[22]) begin
          freeList_22 <= io_retire_prfIdx_1;
        end
        if(_zz_2[23]) begin
          freeList_23 <= io_retire_prfIdx_1;
        end
        if(_zz_2[24]) begin
          freeList_24 <= io_retire_prfIdx_1;
        end
        if(_zz_2[25]) begin
          freeList_25 <= io_retire_prfIdx_1;
        end
        if(_zz_2[26]) begin
          freeList_26 <= io_retire_prfIdx_1;
        end
        if(_zz_2[27]) begin
          freeList_27 <= io_retire_prfIdx_1;
        end
        if(_zz_2[28]) begin
          freeList_28 <= io_retire_prfIdx_1;
        end
        if(_zz_2[29]) begin
          freeList_29 <= io_retire_prfIdx_1;
        end
        if(_zz_2[30]) begin
          freeList_30 <= io_retire_prfIdx_1;
        end
        if(_zz_2[31]) begin
          freeList_31 <= io_retire_prfIdx_1;
        end
        if(_zz_2[32]) begin
          freeList_32 <= io_retire_prfIdx_1;
        end
        if(_zz_2[33]) begin
          freeList_33 <= io_retire_prfIdx_1;
        end
        if(_zz_2[34]) begin
          freeList_34 <= io_retire_prfIdx_1;
        end
        if(_zz_2[35]) begin
          freeList_35 <= io_retire_prfIdx_1;
        end
        if(_zz_2[36]) begin
          freeList_36 <= io_retire_prfIdx_1;
        end
        if(_zz_2[37]) begin
          freeList_37 <= io_retire_prfIdx_1;
        end
        if(_zz_2[38]) begin
          freeList_38 <= io_retire_prfIdx_1;
        end
        if(_zz_2[39]) begin
          freeList_39 <= io_retire_prfIdx_1;
        end
        if(_zz_2[40]) begin
          freeList_40 <= io_retire_prfIdx_1;
        end
        if(_zz_2[41]) begin
          freeList_41 <= io_retire_prfIdx_1;
        end
        if(_zz_2[42]) begin
          freeList_42 <= io_retire_prfIdx_1;
        end
        if(_zz_2[43]) begin
          freeList_43 <= io_retire_prfIdx_1;
        end
        if(_zz_2[44]) begin
          freeList_44 <= io_retire_prfIdx_1;
        end
        if(_zz_2[45]) begin
          freeList_45 <= io_retire_prfIdx_1;
        end
        if(_zz_2[46]) begin
          freeList_46 <= io_retire_prfIdx_1;
        end
        if(_zz_2[47]) begin
          freeList_47 <= io_retire_prfIdx_1;
        end
        if(_zz_2[48]) begin
          freeList_48 <= io_retire_prfIdx_1;
        end
        if(_zz_2[49]) begin
          freeList_49 <= io_retire_prfIdx_1;
        end
        if(_zz_2[50]) begin
          freeList_50 <= io_retire_prfIdx_1;
        end
        if(_zz_2[51]) begin
          freeList_51 <= io_retire_prfIdx_1;
        end
        if(_zz_2[52]) begin
          freeList_52 <= io_retire_prfIdx_1;
        end
        if(_zz_2[53]) begin
          freeList_53 <= io_retire_prfIdx_1;
        end
        if(_zz_2[54]) begin
          freeList_54 <= io_retire_prfIdx_1;
        end
        if(_zz_2[55]) begin
          freeList_55 <= io_retire_prfIdx_1;
        end
        if(_zz_2[56]) begin
          freeList_56 <= io_retire_prfIdx_1;
        end
        if(_zz_2[57]) begin
          freeList_57 <= io_retire_prfIdx_1;
        end
        if(_zz_2[58]) begin
          freeList_58 <= io_retire_prfIdx_1;
        end
        if(_zz_2[59]) begin
          freeList_59 <= io_retire_prfIdx_1;
        end
        if(_zz_2[60]) begin
          freeList_60 <= io_retire_prfIdx_1;
        end
        if(_zz_2[61]) begin
          freeList_61 <= io_retire_prfIdx_1;
        end
        if(_zz_2[62]) begin
          freeList_62 <= io_retire_prfIdx_1;
        end
        if(_zz_2[63]) begin
          freeList_63 <= io_retire_prfIdx_1;
        end
      end
      freePtr_1 <= (freePtr_1 + _zz_freePtr_1);
      retirePtr <= (retirePtr + _zz_retirePtr_1);
      if(io_retire_delayedFlush) begin
        allocPtr_0 <= (retirePtr + 6'h00);
        allocPtr_1 <= (retirePtr + 6'h01);
      end
    end
  end


endmodule

module ARAT (
  input  wire [4:0]    io_retirePort_0_ard,
  input  wire [5:0]    io_retirePort_0_prd,
  input  wire          io_retirePort_0_wen,
  input  wire [4:0]    io_retirePort_1_ard,
  input  wire [5:0]    io_retirePort_1_prd,
  input  wire          io_retirePort_1_wen,
  output wire [5:0]    io_recoveryPort_0,
  output wire [5:0]    io_recoveryPort_1,
  output wire [5:0]    io_recoveryPort_2,
  output wire [5:0]    io_recoveryPort_3,
  output wire [5:0]    io_recoveryPort_4,
  output wire [5:0]    io_recoveryPort_5,
  output wire [5:0]    io_recoveryPort_6,
  output wire [5:0]    io_recoveryPort_7,
  output wire [5:0]    io_recoveryPort_8,
  output wire [5:0]    io_recoveryPort_9,
  output wire [5:0]    io_recoveryPort_10,
  output wire [5:0]    io_recoveryPort_11,
  output wire [5:0]    io_recoveryPort_12,
  output wire [5:0]    io_recoveryPort_13,
  output wire [5:0]    io_recoveryPort_14,
  output wire [5:0]    io_recoveryPort_15,
  output wire [5:0]    io_recoveryPort_16,
  output wire [5:0]    io_recoveryPort_17,
  output wire [5:0]    io_recoveryPort_18,
  output wire [5:0]    io_recoveryPort_19,
  output wire [5:0]    io_recoveryPort_20,
  output wire [5:0]    io_recoveryPort_21,
  output wire [5:0]    io_recoveryPort_22,
  output wire [5:0]    io_recoveryPort_23,
  output wire [5:0]    io_recoveryPort_24,
  output wire [5:0]    io_recoveryPort_25,
  output wire [5:0]    io_recoveryPort_26,
  output wire [5:0]    io_recoveryPort_27,
  output wire [5:0]    io_recoveryPort_28,
  output wire [5:0]    io_recoveryPort_29,
  output wire [5:0]    io_recoveryPort_30,
  output wire [5:0]    io_recoveryPort_31,
  input  wire          aclk,
  input  wire          aresetn
);

  wire       [0:0]    _zz_rat_0;
  wire       [0:0]    _zz_rat_1;
  wire       [0:0]    _zz_rat_2;
  wire       [0:0]    _zz_rat_3;
  wire       [0:0]    _zz_rat_4;
  wire       [0:0]    _zz_rat_5;
  wire       [0:0]    _zz_rat_6;
  wire       [0:0]    _zz_rat_7;
  wire       [0:0]    _zz_rat_8;
  wire       [0:0]    _zz_rat_9;
  wire       [0:0]    _zz_rat_10;
  wire       [0:0]    _zz_rat_11;
  wire       [0:0]    _zz_rat_12;
  wire       [0:0]    _zz_rat_13;
  wire       [0:0]    _zz_rat_14;
  wire       [0:0]    _zz_rat_15;
  wire       [0:0]    _zz_rat_16;
  wire       [0:0]    _zz_rat_17;
  wire       [0:0]    _zz_rat_18;
  wire       [0:0]    _zz_rat_19;
  wire       [0:0]    _zz_rat_20;
  wire       [0:0]    _zz_rat_21;
  wire       [0:0]    _zz_rat_22;
  wire       [0:0]    _zz_rat_23;
  wire       [0:0]    _zz_rat_24;
  wire       [0:0]    _zz_rat_25;
  wire       [0:0]    _zz_rat_26;
  wire       [0:0]    _zz_rat_27;
  wire       [0:0]    _zz_rat_28;
  wire       [0:0]    _zz_rat_29;
  wire       [0:0]    _zz_rat_30;
  wire       [0:0]    _zz_rat_31;
  reg        [5:0]    rat_0;
  reg        [5:0]    rat_1;
  reg        [5:0]    rat_2;
  reg        [5:0]    rat_3;
  reg        [5:0]    rat_4;
  reg        [5:0]    rat_5;
  reg        [5:0]    rat_6;
  reg        [5:0]    rat_7;
  reg        [5:0]    rat_8;
  reg        [5:0]    rat_9;
  reg        [5:0]    rat_10;
  reg        [5:0]    rat_11;
  reg        [5:0]    rat_12;
  reg        [5:0]    rat_13;
  reg        [5:0]    rat_14;
  reg        [5:0]    rat_15;
  reg        [5:0]    rat_16;
  reg        [5:0]    rat_17;
  reg        [5:0]    rat_18;
  reg        [5:0]    rat_19;
  reg        [5:0]    rat_20;
  reg        [5:0]    rat_21;
  reg        [5:0]    rat_22;
  reg        [5:0]    rat_23;
  reg        [5:0]    rat_24;
  reg        [5:0]    rat_25;
  reg        [5:0]    rat_26;
  reg        [5:0]    rat_27;
  reg        [5:0]    rat_28;
  reg        [5:0]    rat_29;
  reg        [5:0]    rat_30;
  reg        [5:0]    rat_31;
  wire       [31:0]   _zz_1;
  wire       [31:0]   _zz_2;

  assign _zz_rat_0 = 1'b0;
  assign _zz_rat_1 = 1'b0;
  assign _zz_rat_2 = 1'b0;
  assign _zz_rat_3 = 1'b0;
  assign _zz_rat_4 = 1'b0;
  assign _zz_rat_5 = 1'b0;
  assign _zz_rat_6 = 1'b0;
  assign _zz_rat_7 = 1'b0;
  assign _zz_rat_8 = 1'b0;
  assign _zz_rat_9 = 1'b0;
  assign _zz_rat_10 = 1'b0;
  assign _zz_rat_11 = 1'b0;
  assign _zz_rat_12 = 1'b0;
  assign _zz_rat_13 = 1'b0;
  assign _zz_rat_14 = 1'b0;
  assign _zz_rat_15 = 1'b0;
  assign _zz_rat_16 = 1'b0;
  assign _zz_rat_17 = 1'b0;
  assign _zz_rat_18 = 1'b0;
  assign _zz_rat_19 = 1'b0;
  assign _zz_rat_20 = 1'b0;
  assign _zz_rat_21 = 1'b0;
  assign _zz_rat_22 = 1'b0;
  assign _zz_rat_23 = 1'b0;
  assign _zz_rat_24 = 1'b0;
  assign _zz_rat_25 = 1'b0;
  assign _zz_rat_26 = 1'b0;
  assign _zz_rat_27 = 1'b0;
  assign _zz_rat_28 = 1'b0;
  assign _zz_rat_29 = 1'b0;
  assign _zz_rat_30 = 1'b0;
  assign _zz_rat_31 = 1'b0;
  assign _zz_1 = ({31'd0,1'b1} <<< io_retirePort_0_ard);
  assign _zz_2 = ({31'd0,1'b1} <<< io_retirePort_1_ard);
  assign io_recoveryPort_0 = rat_0;
  assign io_recoveryPort_1 = rat_1;
  assign io_recoveryPort_2 = rat_2;
  assign io_recoveryPort_3 = rat_3;
  assign io_recoveryPort_4 = rat_4;
  assign io_recoveryPort_5 = rat_5;
  assign io_recoveryPort_6 = rat_6;
  assign io_recoveryPort_7 = rat_7;
  assign io_recoveryPort_8 = rat_8;
  assign io_recoveryPort_9 = rat_9;
  assign io_recoveryPort_10 = rat_10;
  assign io_recoveryPort_11 = rat_11;
  assign io_recoveryPort_12 = rat_12;
  assign io_recoveryPort_13 = rat_13;
  assign io_recoveryPort_14 = rat_14;
  assign io_recoveryPort_15 = rat_15;
  assign io_recoveryPort_16 = rat_16;
  assign io_recoveryPort_17 = rat_17;
  assign io_recoveryPort_18 = rat_18;
  assign io_recoveryPort_19 = rat_19;
  assign io_recoveryPort_20 = rat_20;
  assign io_recoveryPort_21 = rat_21;
  assign io_recoveryPort_22 = rat_22;
  assign io_recoveryPort_23 = rat_23;
  assign io_recoveryPort_24 = rat_24;
  assign io_recoveryPort_25 = rat_25;
  assign io_recoveryPort_26 = rat_26;
  assign io_recoveryPort_27 = rat_27;
  assign io_recoveryPort_28 = rat_28;
  assign io_recoveryPort_29 = rat_29;
  assign io_recoveryPort_30 = rat_30;
  assign io_recoveryPort_31 = rat_31;
  always @(posedge aclk) begin
    if(!aresetn) begin
      rat_0 <= {5'd0, _zz_rat_0};
      rat_1 <= {5'd0, _zz_rat_1};
      rat_2 <= {5'd0, _zz_rat_2};
      rat_3 <= {5'd0, _zz_rat_3};
      rat_4 <= {5'd0, _zz_rat_4};
      rat_5 <= {5'd0, _zz_rat_5};
      rat_6 <= {5'd0, _zz_rat_6};
      rat_7 <= {5'd0, _zz_rat_7};
      rat_8 <= {5'd0, _zz_rat_8};
      rat_9 <= {5'd0, _zz_rat_9};
      rat_10 <= {5'd0, _zz_rat_10};
      rat_11 <= {5'd0, _zz_rat_11};
      rat_12 <= {5'd0, _zz_rat_12};
      rat_13 <= {5'd0, _zz_rat_13};
      rat_14 <= {5'd0, _zz_rat_14};
      rat_15 <= {5'd0, _zz_rat_15};
      rat_16 <= {5'd0, _zz_rat_16};
      rat_17 <= {5'd0, _zz_rat_17};
      rat_18 <= {5'd0, _zz_rat_18};
      rat_19 <= {5'd0, _zz_rat_19};
      rat_20 <= {5'd0, _zz_rat_20};
      rat_21 <= {5'd0, _zz_rat_21};
      rat_22 <= {5'd0, _zz_rat_22};
      rat_23 <= {5'd0, _zz_rat_23};
      rat_24 <= {5'd0, _zz_rat_24};
      rat_25 <= {5'd0, _zz_rat_25};
      rat_26 <= {5'd0, _zz_rat_26};
      rat_27 <= {5'd0, _zz_rat_27};
      rat_28 <= {5'd0, _zz_rat_28};
      rat_29 <= {5'd0, _zz_rat_29};
      rat_30 <= {5'd0, _zz_rat_30};
      rat_31 <= {5'd0, _zz_rat_31};
    end else begin
      if(io_retirePort_0_wen) begin
        if(_zz_1[0]) begin
          rat_0 <= io_retirePort_0_prd;
        end
        if(_zz_1[1]) begin
          rat_1 <= io_retirePort_0_prd;
        end
        if(_zz_1[2]) begin
          rat_2 <= io_retirePort_0_prd;
        end
        if(_zz_1[3]) begin
          rat_3 <= io_retirePort_0_prd;
        end
        if(_zz_1[4]) begin
          rat_4 <= io_retirePort_0_prd;
        end
        if(_zz_1[5]) begin
          rat_5 <= io_retirePort_0_prd;
        end
        if(_zz_1[6]) begin
          rat_6 <= io_retirePort_0_prd;
        end
        if(_zz_1[7]) begin
          rat_7 <= io_retirePort_0_prd;
        end
        if(_zz_1[8]) begin
          rat_8 <= io_retirePort_0_prd;
        end
        if(_zz_1[9]) begin
          rat_9 <= io_retirePort_0_prd;
        end
        if(_zz_1[10]) begin
          rat_10 <= io_retirePort_0_prd;
        end
        if(_zz_1[11]) begin
          rat_11 <= io_retirePort_0_prd;
        end
        if(_zz_1[12]) begin
          rat_12 <= io_retirePort_0_prd;
        end
        if(_zz_1[13]) begin
          rat_13 <= io_retirePort_0_prd;
        end
        if(_zz_1[14]) begin
          rat_14 <= io_retirePort_0_prd;
        end
        if(_zz_1[15]) begin
          rat_15 <= io_retirePort_0_prd;
        end
        if(_zz_1[16]) begin
          rat_16 <= io_retirePort_0_prd;
        end
        if(_zz_1[17]) begin
          rat_17 <= io_retirePort_0_prd;
        end
        if(_zz_1[18]) begin
          rat_18 <= io_retirePort_0_prd;
        end
        if(_zz_1[19]) begin
          rat_19 <= io_retirePort_0_prd;
        end
        if(_zz_1[20]) begin
          rat_20 <= io_retirePort_0_prd;
        end
        if(_zz_1[21]) begin
          rat_21 <= io_retirePort_0_prd;
        end
        if(_zz_1[22]) begin
          rat_22 <= io_retirePort_0_prd;
        end
        if(_zz_1[23]) begin
          rat_23 <= io_retirePort_0_prd;
        end
        if(_zz_1[24]) begin
          rat_24 <= io_retirePort_0_prd;
        end
        if(_zz_1[25]) begin
          rat_25 <= io_retirePort_0_prd;
        end
        if(_zz_1[26]) begin
          rat_26 <= io_retirePort_0_prd;
        end
        if(_zz_1[27]) begin
          rat_27 <= io_retirePort_0_prd;
        end
        if(_zz_1[28]) begin
          rat_28 <= io_retirePort_0_prd;
        end
        if(_zz_1[29]) begin
          rat_29 <= io_retirePort_0_prd;
        end
        if(_zz_1[30]) begin
          rat_30 <= io_retirePort_0_prd;
        end
        if(_zz_1[31]) begin
          rat_31 <= io_retirePort_0_prd;
        end
      end
      if(io_retirePort_1_wen) begin
        if(_zz_2[0]) begin
          rat_0 <= io_retirePort_1_prd;
        end
        if(_zz_2[1]) begin
          rat_1 <= io_retirePort_1_prd;
        end
        if(_zz_2[2]) begin
          rat_2 <= io_retirePort_1_prd;
        end
        if(_zz_2[3]) begin
          rat_3 <= io_retirePort_1_prd;
        end
        if(_zz_2[4]) begin
          rat_4 <= io_retirePort_1_prd;
        end
        if(_zz_2[5]) begin
          rat_5 <= io_retirePort_1_prd;
        end
        if(_zz_2[6]) begin
          rat_6 <= io_retirePort_1_prd;
        end
        if(_zz_2[7]) begin
          rat_7 <= io_retirePort_1_prd;
        end
        if(_zz_2[8]) begin
          rat_8 <= io_retirePort_1_prd;
        end
        if(_zz_2[9]) begin
          rat_9 <= io_retirePort_1_prd;
        end
        if(_zz_2[10]) begin
          rat_10 <= io_retirePort_1_prd;
        end
        if(_zz_2[11]) begin
          rat_11 <= io_retirePort_1_prd;
        end
        if(_zz_2[12]) begin
          rat_12 <= io_retirePort_1_prd;
        end
        if(_zz_2[13]) begin
          rat_13 <= io_retirePort_1_prd;
        end
        if(_zz_2[14]) begin
          rat_14 <= io_retirePort_1_prd;
        end
        if(_zz_2[15]) begin
          rat_15 <= io_retirePort_1_prd;
        end
        if(_zz_2[16]) begin
          rat_16 <= io_retirePort_1_prd;
        end
        if(_zz_2[17]) begin
          rat_17 <= io_retirePort_1_prd;
        end
        if(_zz_2[18]) begin
          rat_18 <= io_retirePort_1_prd;
        end
        if(_zz_2[19]) begin
          rat_19 <= io_retirePort_1_prd;
        end
        if(_zz_2[20]) begin
          rat_20 <= io_retirePort_1_prd;
        end
        if(_zz_2[21]) begin
          rat_21 <= io_retirePort_1_prd;
        end
        if(_zz_2[22]) begin
          rat_22 <= io_retirePort_1_prd;
        end
        if(_zz_2[23]) begin
          rat_23 <= io_retirePort_1_prd;
        end
        if(_zz_2[24]) begin
          rat_24 <= io_retirePort_1_prd;
        end
        if(_zz_2[25]) begin
          rat_25 <= io_retirePort_1_prd;
        end
        if(_zz_2[26]) begin
          rat_26 <= io_retirePort_1_prd;
        end
        if(_zz_2[27]) begin
          rat_27 <= io_retirePort_1_prd;
        end
        if(_zz_2[28]) begin
          rat_28 <= io_retirePort_1_prd;
        end
        if(_zz_2[29]) begin
          rat_29 <= io_retirePort_1_prd;
        end
        if(_zz_2[30]) begin
          rat_30 <= io_retirePort_1_prd;
        end
        if(_zz_2[31]) begin
          rat_31 <= io_retirePort_1_prd;
        end
      end
    end
  end


endmodule

module SRAT (
  input  wire [4:0]    io_writePort_0_ard,
  input  wire [5:0]    io_writePort_0_prd,
  input  wire          io_writePort_0_wen,
  input  wire [4:0]    io_writePort_1_ard,
  input  wire [5:0]    io_writePort_1_prd,
  input  wire          io_writePort_1_wen,
  input  wire [5:0]    io_updatePort_0_prd,
  input  wire          io_updatePort_0_wen,
  input  wire [5:0]    io_updatePort_1_prd,
  input  wire          io_updatePort_1_wen,
  input  wire [5:0]    io_updatePort_2_prd,
  input  wire          io_updatePort_2_wen,
  input  wire [5:0]    io_updatePort_3_prd,
  input  wire          io_updatePort_3_wen,
  input  wire [5:0]    io_updatePort_4_prd,
  input  wire          io_updatePort_4_wen,
  input  wire [4:0]    io_srcReadPort_0_0_ard,
  output wire [5:0]    io_srcReadPort_0_0_prd,
  output wire          io_srcReadPort_0_0_valid,
  input  wire [4:0]    io_srcReadPort_0_1_ard,
  output wire [5:0]    io_srcReadPort_0_1_prd,
  output wire          io_srcReadPort_0_1_valid,
  input  wire [4:0]    io_srcReadPort_1_0_ard,
  output wire [5:0]    io_srcReadPort_1_0_prd,
  output wire          io_srcReadPort_1_0_valid,
  input  wire [4:0]    io_srcReadPort_1_1_ard,
  output wire [5:0]    io_srcReadPort_1_1_prd,
  output wire          io_srcReadPort_1_1_valid,
  input  wire [4:0]    io_prevPRDReadPort_0_ard,
  output wire [5:0]    io_prevPRDReadPort_0_prd,
  output wire          io_prevPRDReadPort_0_valid,
  input  wire [4:0]    io_prevPRDReadPort_1_ard,
  output wire [5:0]    io_prevPRDReadPort_1_prd,
  output wire          io_prevPRDReadPort_1_valid,
  input  wire          io_delayedRecovery,
  input  wire [5:0]    io_recoveryPort_0,
  input  wire [5:0]    io_recoveryPort_1,
  input  wire [5:0]    io_recoveryPort_2,
  input  wire [5:0]    io_recoveryPort_3,
  input  wire [5:0]    io_recoveryPort_4,
  input  wire [5:0]    io_recoveryPort_5,
  input  wire [5:0]    io_recoveryPort_6,
  input  wire [5:0]    io_recoveryPort_7,
  input  wire [5:0]    io_recoveryPort_8,
  input  wire [5:0]    io_recoveryPort_9,
  input  wire [5:0]    io_recoveryPort_10,
  input  wire [5:0]    io_recoveryPort_11,
  input  wire [5:0]    io_recoveryPort_12,
  input  wire [5:0]    io_recoveryPort_13,
  input  wire [5:0]    io_recoveryPort_14,
  input  wire [5:0]    io_recoveryPort_15,
  input  wire [5:0]    io_recoveryPort_16,
  input  wire [5:0]    io_recoveryPort_17,
  input  wire [5:0]    io_recoveryPort_18,
  input  wire [5:0]    io_recoveryPort_19,
  input  wire [5:0]    io_recoveryPort_20,
  input  wire [5:0]    io_recoveryPort_21,
  input  wire [5:0]    io_recoveryPort_22,
  input  wire [5:0]    io_recoveryPort_23,
  input  wire [5:0]    io_recoveryPort_24,
  input  wire [5:0]    io_recoveryPort_25,
  input  wire [5:0]    io_recoveryPort_26,
  input  wire [5:0]    io_recoveryPort_27,
  input  wire [5:0]    io_recoveryPort_28,
  input  wire [5:0]    io_recoveryPort_29,
  input  wire [5:0]    io_recoveryPort_30,
  input  wire [5:0]    io_recoveryPort_31,
  input  wire          aclk,
  input  wire          aresetn
);

  wire       [0:0]    _zz_rat_0_prfIdx;
  wire       [0:0]    _zz_rat_1_prfIdx;
  wire       [0:0]    _zz_rat_2_prfIdx;
  wire       [0:0]    _zz_rat_3_prfIdx;
  wire       [0:0]    _zz_rat_4_prfIdx;
  wire       [0:0]    _zz_rat_5_prfIdx;
  wire       [0:0]    _zz_rat_6_prfIdx;
  wire       [0:0]    _zz_rat_7_prfIdx;
  wire       [0:0]    _zz_rat_8_prfIdx;
  wire       [0:0]    _zz_rat_9_prfIdx;
  wire       [0:0]    _zz_rat_10_prfIdx;
  wire       [0:0]    _zz_rat_11_prfIdx;
  wire       [0:0]    _zz_rat_12_prfIdx;
  wire       [0:0]    _zz_rat_13_prfIdx;
  wire       [0:0]    _zz_rat_14_prfIdx;
  wire       [0:0]    _zz_rat_15_prfIdx;
  wire       [0:0]    _zz_rat_16_prfIdx;
  wire       [0:0]    _zz_rat_17_prfIdx;
  wire       [0:0]    _zz_rat_18_prfIdx;
  wire       [0:0]    _zz_rat_19_prfIdx;
  wire       [0:0]    _zz_rat_20_prfIdx;
  wire       [0:0]    _zz_rat_21_prfIdx;
  wire       [0:0]    _zz_rat_22_prfIdx;
  wire       [0:0]    _zz_rat_23_prfIdx;
  wire       [0:0]    _zz_rat_24_prfIdx;
  wire       [0:0]    _zz_rat_25_prfIdx;
  wire       [0:0]    _zz_rat_26_prfIdx;
  wire       [0:0]    _zz_rat_27_prfIdx;
  wire       [0:0]    _zz_rat_28_prfIdx;
  wire       [0:0]    _zz_rat_29_prfIdx;
  wire       [0:0]    _zz_rat_30_prfIdx;
  wire       [0:0]    _zz_rat_31_prfIdx;
  reg        [5:0]    _zz_io_srcReadPort_0_0_prd;
  wire       [4:0]    _zz_io_srcReadPort_0_0_prd_1;
  reg                 _zz_io_srcReadPort_0_0_valid;
  wire       [4:0]    _zz_io_srcReadPort_0_0_valid_1;
  reg        [5:0]    _zz_io_srcReadPort_0_1_prd;
  wire       [4:0]    _zz_io_srcReadPort_0_1_prd_1;
  reg                 _zz_io_srcReadPort_0_1_valid;
  wire       [4:0]    _zz_io_srcReadPort_0_1_valid_1;
  reg        [5:0]    _zz_io_srcReadPort_1_0_prd;
  wire       [4:0]    _zz_io_srcReadPort_1_0_prd_1;
  reg                 _zz_io_srcReadPort_1_0_valid;
  wire       [4:0]    _zz_io_srcReadPort_1_0_valid_1;
  reg        [5:0]    _zz_io_srcReadPort_1_1_prd;
  wire       [4:0]    _zz_io_srcReadPort_1_1_prd_1;
  reg                 _zz_io_srcReadPort_1_1_valid;
  wire       [4:0]    _zz_io_srcReadPort_1_1_valid_1;
  reg        [5:0]    _zz_io_prevPRDReadPort_0_prd;
  wire       [4:0]    _zz_io_prevPRDReadPort_0_prd_1;
  reg                 _zz_io_prevPRDReadPort_0_valid;
  wire       [4:0]    _zz_io_prevPRDReadPort_0_valid_1;
  reg        [5:0]    _zz_io_prevPRDReadPort_1_prd;
  wire       [4:0]    _zz_io_prevPRDReadPort_1_prd_1;
  reg                 _zz_io_prevPRDReadPort_1_valid;
  wire       [4:0]    _zz_io_prevPRDReadPort_1_valid_1;
  reg        [5:0]    rat_0_prfIdx;
  reg                 rat_0_valid;
  reg        [5:0]    rat_1_prfIdx;
  reg                 rat_1_valid;
  reg        [5:0]    rat_2_prfIdx;
  reg                 rat_2_valid;
  reg        [5:0]    rat_3_prfIdx;
  reg                 rat_3_valid;
  reg        [5:0]    rat_4_prfIdx;
  reg                 rat_4_valid;
  reg        [5:0]    rat_5_prfIdx;
  reg                 rat_5_valid;
  reg        [5:0]    rat_6_prfIdx;
  reg                 rat_6_valid;
  reg        [5:0]    rat_7_prfIdx;
  reg                 rat_7_valid;
  reg        [5:0]    rat_8_prfIdx;
  reg                 rat_8_valid;
  reg        [5:0]    rat_9_prfIdx;
  reg                 rat_9_valid;
  reg        [5:0]    rat_10_prfIdx;
  reg                 rat_10_valid;
  reg        [5:0]    rat_11_prfIdx;
  reg                 rat_11_valid;
  reg        [5:0]    rat_12_prfIdx;
  reg                 rat_12_valid;
  reg        [5:0]    rat_13_prfIdx;
  reg                 rat_13_valid;
  reg        [5:0]    rat_14_prfIdx;
  reg                 rat_14_valid;
  reg        [5:0]    rat_15_prfIdx;
  reg                 rat_15_valid;
  reg        [5:0]    rat_16_prfIdx;
  reg                 rat_16_valid;
  reg        [5:0]    rat_17_prfIdx;
  reg                 rat_17_valid;
  reg        [5:0]    rat_18_prfIdx;
  reg                 rat_18_valid;
  reg        [5:0]    rat_19_prfIdx;
  reg                 rat_19_valid;
  reg        [5:0]    rat_20_prfIdx;
  reg                 rat_20_valid;
  reg        [5:0]    rat_21_prfIdx;
  reg                 rat_21_valid;
  reg        [5:0]    rat_22_prfIdx;
  reg                 rat_22_valid;
  reg        [5:0]    rat_23_prfIdx;
  reg                 rat_23_valid;
  reg        [5:0]    rat_24_prfIdx;
  reg                 rat_24_valid;
  reg        [5:0]    rat_25_prfIdx;
  reg                 rat_25_valid;
  reg        [5:0]    rat_26_prfIdx;
  reg                 rat_26_valid;
  reg        [5:0]    rat_27_prfIdx;
  reg                 rat_27_valid;
  reg        [5:0]    rat_28_prfIdx;
  reg                 rat_28_valid;
  reg        [5:0]    rat_29_prfIdx;
  reg                 rat_29_valid;
  reg        [5:0]    rat_30_prfIdx;
  reg                 rat_30_valid;
  reg        [5:0]    rat_31_prfIdx;
  reg                 rat_31_valid;
  wire                when_RAT_l30;
  wire                when_RAT_l30_1;
  wire                when_RAT_l30_2;
  wire                when_RAT_l30_3;
  wire                when_RAT_l30_4;
  wire                when_RAT_l30_5;
  wire                when_RAT_l30_6;
  wire                when_RAT_l30_7;
  wire                when_RAT_l30_8;
  wire                when_RAT_l30_9;
  wire                when_RAT_l30_10;
  wire                when_RAT_l30_11;
  wire                when_RAT_l30_12;
  wire                when_RAT_l30_13;
  wire                when_RAT_l30_14;
  wire                when_RAT_l30_15;
  wire                when_RAT_l30_16;
  wire                when_RAT_l30_17;
  wire                when_RAT_l30_18;
  wire                when_RAT_l30_19;
  wire                when_RAT_l30_20;
  wire                when_RAT_l30_21;
  wire                when_RAT_l30_22;
  wire                when_RAT_l30_23;
  wire                when_RAT_l30_24;
  wire                when_RAT_l30_25;
  wire                when_RAT_l30_26;
  wire                when_RAT_l30_27;
  wire                when_RAT_l30_28;
  wire                when_RAT_l30_29;
  wire                when_RAT_l30_30;
  wire                when_RAT_l30_31;
  wire                when_RAT_l30_32;
  wire                when_RAT_l30_33;
  wire                when_RAT_l30_34;
  wire                when_RAT_l30_35;
  wire                when_RAT_l30_36;
  wire                when_RAT_l30_37;
  wire                when_RAT_l30_38;
  wire                when_RAT_l30_39;
  wire                when_RAT_l30_40;
  wire                when_RAT_l30_41;
  wire                when_RAT_l30_42;
  wire                when_RAT_l30_43;
  wire                when_RAT_l30_44;
  wire                when_RAT_l30_45;
  wire                when_RAT_l30_46;
  wire                when_RAT_l30_47;
  wire                when_RAT_l30_48;
  wire                when_RAT_l30_49;
  wire                when_RAT_l30_50;
  wire                when_RAT_l30_51;
  wire                when_RAT_l30_52;
  wire                when_RAT_l30_53;
  wire                when_RAT_l30_54;
  wire                when_RAT_l30_55;
  wire                when_RAT_l30_56;
  wire                when_RAT_l30_57;
  wire                when_RAT_l30_58;
  wire                when_RAT_l30_59;
  wire                when_RAT_l30_60;
  wire                when_RAT_l30_61;
  wire                when_RAT_l30_62;
  wire                when_RAT_l30_63;
  wire                when_RAT_l30_64;
  wire                when_RAT_l30_65;
  wire                when_RAT_l30_66;
  wire                when_RAT_l30_67;
  wire                when_RAT_l30_68;
  wire                when_RAT_l30_69;
  wire                when_RAT_l30_70;
  wire                when_RAT_l30_71;
  wire                when_RAT_l30_72;
  wire                when_RAT_l30_73;
  wire                when_RAT_l30_74;
  wire                when_RAT_l30_75;
  wire                when_RAT_l30_76;
  wire                when_RAT_l30_77;
  wire                when_RAT_l30_78;
  wire                when_RAT_l30_79;
  wire                when_RAT_l30_80;
  wire                when_RAT_l30_81;
  wire                when_RAT_l30_82;
  wire                when_RAT_l30_83;
  wire                when_RAT_l30_84;
  wire                when_RAT_l30_85;
  wire                when_RAT_l30_86;
  wire                when_RAT_l30_87;
  wire                when_RAT_l30_88;
  wire                when_RAT_l30_89;
  wire                when_RAT_l30_90;
  wire                when_RAT_l30_91;
  wire                when_RAT_l30_92;
  wire                when_RAT_l30_93;
  wire                when_RAT_l30_94;
  wire                when_RAT_l30_95;
  wire                when_RAT_l30_96;
  wire                when_RAT_l30_97;
  wire                when_RAT_l30_98;
  wire                when_RAT_l30_99;
  wire                when_RAT_l30_100;
  wire                when_RAT_l30_101;
  wire                when_RAT_l30_102;
  wire                when_RAT_l30_103;
  wire                when_RAT_l30_104;
  wire                when_RAT_l30_105;
  wire                when_RAT_l30_106;
  wire                when_RAT_l30_107;
  wire                when_RAT_l30_108;
  wire                when_RAT_l30_109;
  wire                when_RAT_l30_110;
  wire                when_RAT_l30_111;
  wire                when_RAT_l30_112;
  wire                when_RAT_l30_113;
  wire                when_RAT_l30_114;
  wire                when_RAT_l30_115;
  wire                when_RAT_l30_116;
  wire                when_RAT_l30_117;
  wire                when_RAT_l30_118;
  wire                when_RAT_l30_119;
  wire                when_RAT_l30_120;
  wire                when_RAT_l30_121;
  wire                when_RAT_l30_122;
  wire                when_RAT_l30_123;
  wire                when_RAT_l30_124;
  wire                when_RAT_l30_125;
  wire                when_RAT_l30_126;
  wire                when_RAT_l30_127;
  wire                when_RAT_l30_128;
  wire                when_RAT_l30_129;
  wire                when_RAT_l30_130;
  wire                when_RAT_l30_131;
  wire                when_RAT_l30_132;
  wire                when_RAT_l30_133;
  wire                when_RAT_l30_134;
  wire                when_RAT_l30_135;
  wire                when_RAT_l30_136;
  wire                when_RAT_l30_137;
  wire                when_RAT_l30_138;
  wire                when_RAT_l30_139;
  wire                when_RAT_l30_140;
  wire                when_RAT_l30_141;
  wire                when_RAT_l30_142;
  wire                when_RAT_l30_143;
  wire                when_RAT_l30_144;
  wire                when_RAT_l30_145;
  wire                when_RAT_l30_146;
  wire                when_RAT_l30_147;
  wire                when_RAT_l30_148;
  wire                when_RAT_l30_149;
  wire                when_RAT_l30_150;
  wire                when_RAT_l30_151;
  wire                when_RAT_l30_152;
  wire                when_RAT_l30_153;
  wire                when_RAT_l30_154;
  wire                when_RAT_l30_155;
  wire                when_RAT_l30_156;
  wire                when_RAT_l30_157;
  wire                when_RAT_l30_158;
  wire                when_RAT_l30_159;
  wire       [31:0]   _zz_1;
  wire       [31:0]   _zz_2;
  wire       [31:0]   _zz_3;
  wire       [31:0]   _zz_4;

  assign _zz_rat_0_prfIdx = 1'b0;
  assign _zz_rat_1_prfIdx = 1'b0;
  assign _zz_rat_2_prfIdx = 1'b0;
  assign _zz_rat_3_prfIdx = 1'b0;
  assign _zz_rat_4_prfIdx = 1'b0;
  assign _zz_rat_5_prfIdx = 1'b0;
  assign _zz_rat_6_prfIdx = 1'b0;
  assign _zz_rat_7_prfIdx = 1'b0;
  assign _zz_rat_8_prfIdx = 1'b0;
  assign _zz_rat_9_prfIdx = 1'b0;
  assign _zz_rat_10_prfIdx = 1'b0;
  assign _zz_rat_11_prfIdx = 1'b0;
  assign _zz_rat_12_prfIdx = 1'b0;
  assign _zz_rat_13_prfIdx = 1'b0;
  assign _zz_rat_14_prfIdx = 1'b0;
  assign _zz_rat_15_prfIdx = 1'b0;
  assign _zz_rat_16_prfIdx = 1'b0;
  assign _zz_rat_17_prfIdx = 1'b0;
  assign _zz_rat_18_prfIdx = 1'b0;
  assign _zz_rat_19_prfIdx = 1'b0;
  assign _zz_rat_20_prfIdx = 1'b0;
  assign _zz_rat_21_prfIdx = 1'b0;
  assign _zz_rat_22_prfIdx = 1'b0;
  assign _zz_rat_23_prfIdx = 1'b0;
  assign _zz_rat_24_prfIdx = 1'b0;
  assign _zz_rat_25_prfIdx = 1'b0;
  assign _zz_rat_26_prfIdx = 1'b0;
  assign _zz_rat_27_prfIdx = 1'b0;
  assign _zz_rat_28_prfIdx = 1'b0;
  assign _zz_rat_29_prfIdx = 1'b0;
  assign _zz_rat_30_prfIdx = 1'b0;
  assign _zz_rat_31_prfIdx = 1'b0;
  assign _zz_io_srcReadPort_0_0_prd_1 = io_srcReadPort_0_0_ard;
  assign _zz_io_srcReadPort_0_0_valid_1 = io_srcReadPort_0_0_ard;
  assign _zz_io_srcReadPort_0_1_prd_1 = io_srcReadPort_0_1_ard;
  assign _zz_io_srcReadPort_0_1_valid_1 = io_srcReadPort_0_1_ard;
  assign _zz_io_srcReadPort_1_0_prd_1 = io_srcReadPort_1_0_ard;
  assign _zz_io_srcReadPort_1_0_valid_1 = io_srcReadPort_1_0_ard;
  assign _zz_io_srcReadPort_1_1_prd_1 = io_srcReadPort_1_1_ard;
  assign _zz_io_srcReadPort_1_1_valid_1 = io_srcReadPort_1_1_ard;
  assign _zz_io_prevPRDReadPort_0_prd_1 = io_prevPRDReadPort_0_ard;
  assign _zz_io_prevPRDReadPort_0_valid_1 = io_prevPRDReadPort_0_ard;
  assign _zz_io_prevPRDReadPort_1_prd_1 = io_prevPRDReadPort_1_ard;
  assign _zz_io_prevPRDReadPort_1_valid_1 = io_prevPRDReadPort_1_ard;
  always @(*) begin
    case(_zz_io_srcReadPort_0_0_prd_1)
      5'b00000 : _zz_io_srcReadPort_0_0_prd = rat_0_prfIdx;
      5'b00001 : _zz_io_srcReadPort_0_0_prd = rat_1_prfIdx;
      5'b00010 : _zz_io_srcReadPort_0_0_prd = rat_2_prfIdx;
      5'b00011 : _zz_io_srcReadPort_0_0_prd = rat_3_prfIdx;
      5'b00100 : _zz_io_srcReadPort_0_0_prd = rat_4_prfIdx;
      5'b00101 : _zz_io_srcReadPort_0_0_prd = rat_5_prfIdx;
      5'b00110 : _zz_io_srcReadPort_0_0_prd = rat_6_prfIdx;
      5'b00111 : _zz_io_srcReadPort_0_0_prd = rat_7_prfIdx;
      5'b01000 : _zz_io_srcReadPort_0_0_prd = rat_8_prfIdx;
      5'b01001 : _zz_io_srcReadPort_0_0_prd = rat_9_prfIdx;
      5'b01010 : _zz_io_srcReadPort_0_0_prd = rat_10_prfIdx;
      5'b01011 : _zz_io_srcReadPort_0_0_prd = rat_11_prfIdx;
      5'b01100 : _zz_io_srcReadPort_0_0_prd = rat_12_prfIdx;
      5'b01101 : _zz_io_srcReadPort_0_0_prd = rat_13_prfIdx;
      5'b01110 : _zz_io_srcReadPort_0_0_prd = rat_14_prfIdx;
      5'b01111 : _zz_io_srcReadPort_0_0_prd = rat_15_prfIdx;
      5'b10000 : _zz_io_srcReadPort_0_0_prd = rat_16_prfIdx;
      5'b10001 : _zz_io_srcReadPort_0_0_prd = rat_17_prfIdx;
      5'b10010 : _zz_io_srcReadPort_0_0_prd = rat_18_prfIdx;
      5'b10011 : _zz_io_srcReadPort_0_0_prd = rat_19_prfIdx;
      5'b10100 : _zz_io_srcReadPort_0_0_prd = rat_20_prfIdx;
      5'b10101 : _zz_io_srcReadPort_0_0_prd = rat_21_prfIdx;
      5'b10110 : _zz_io_srcReadPort_0_0_prd = rat_22_prfIdx;
      5'b10111 : _zz_io_srcReadPort_0_0_prd = rat_23_prfIdx;
      5'b11000 : _zz_io_srcReadPort_0_0_prd = rat_24_prfIdx;
      5'b11001 : _zz_io_srcReadPort_0_0_prd = rat_25_prfIdx;
      5'b11010 : _zz_io_srcReadPort_0_0_prd = rat_26_prfIdx;
      5'b11011 : _zz_io_srcReadPort_0_0_prd = rat_27_prfIdx;
      5'b11100 : _zz_io_srcReadPort_0_0_prd = rat_28_prfIdx;
      5'b11101 : _zz_io_srcReadPort_0_0_prd = rat_29_prfIdx;
      5'b11110 : _zz_io_srcReadPort_0_0_prd = rat_30_prfIdx;
      default : _zz_io_srcReadPort_0_0_prd = rat_31_prfIdx;
    endcase
  end

  always @(*) begin
    case(_zz_io_srcReadPort_0_0_valid_1)
      5'b00000 : _zz_io_srcReadPort_0_0_valid = rat_0_valid;
      5'b00001 : _zz_io_srcReadPort_0_0_valid = rat_1_valid;
      5'b00010 : _zz_io_srcReadPort_0_0_valid = rat_2_valid;
      5'b00011 : _zz_io_srcReadPort_0_0_valid = rat_3_valid;
      5'b00100 : _zz_io_srcReadPort_0_0_valid = rat_4_valid;
      5'b00101 : _zz_io_srcReadPort_0_0_valid = rat_5_valid;
      5'b00110 : _zz_io_srcReadPort_0_0_valid = rat_6_valid;
      5'b00111 : _zz_io_srcReadPort_0_0_valid = rat_7_valid;
      5'b01000 : _zz_io_srcReadPort_0_0_valid = rat_8_valid;
      5'b01001 : _zz_io_srcReadPort_0_0_valid = rat_9_valid;
      5'b01010 : _zz_io_srcReadPort_0_0_valid = rat_10_valid;
      5'b01011 : _zz_io_srcReadPort_0_0_valid = rat_11_valid;
      5'b01100 : _zz_io_srcReadPort_0_0_valid = rat_12_valid;
      5'b01101 : _zz_io_srcReadPort_0_0_valid = rat_13_valid;
      5'b01110 : _zz_io_srcReadPort_0_0_valid = rat_14_valid;
      5'b01111 : _zz_io_srcReadPort_0_0_valid = rat_15_valid;
      5'b10000 : _zz_io_srcReadPort_0_0_valid = rat_16_valid;
      5'b10001 : _zz_io_srcReadPort_0_0_valid = rat_17_valid;
      5'b10010 : _zz_io_srcReadPort_0_0_valid = rat_18_valid;
      5'b10011 : _zz_io_srcReadPort_0_0_valid = rat_19_valid;
      5'b10100 : _zz_io_srcReadPort_0_0_valid = rat_20_valid;
      5'b10101 : _zz_io_srcReadPort_0_0_valid = rat_21_valid;
      5'b10110 : _zz_io_srcReadPort_0_0_valid = rat_22_valid;
      5'b10111 : _zz_io_srcReadPort_0_0_valid = rat_23_valid;
      5'b11000 : _zz_io_srcReadPort_0_0_valid = rat_24_valid;
      5'b11001 : _zz_io_srcReadPort_0_0_valid = rat_25_valid;
      5'b11010 : _zz_io_srcReadPort_0_0_valid = rat_26_valid;
      5'b11011 : _zz_io_srcReadPort_0_0_valid = rat_27_valid;
      5'b11100 : _zz_io_srcReadPort_0_0_valid = rat_28_valid;
      5'b11101 : _zz_io_srcReadPort_0_0_valid = rat_29_valid;
      5'b11110 : _zz_io_srcReadPort_0_0_valid = rat_30_valid;
      default : _zz_io_srcReadPort_0_0_valid = rat_31_valid;
    endcase
  end

  always @(*) begin
    case(_zz_io_srcReadPort_0_1_prd_1)
      5'b00000 : _zz_io_srcReadPort_0_1_prd = rat_0_prfIdx;
      5'b00001 : _zz_io_srcReadPort_0_1_prd = rat_1_prfIdx;
      5'b00010 : _zz_io_srcReadPort_0_1_prd = rat_2_prfIdx;
      5'b00011 : _zz_io_srcReadPort_0_1_prd = rat_3_prfIdx;
      5'b00100 : _zz_io_srcReadPort_0_1_prd = rat_4_prfIdx;
      5'b00101 : _zz_io_srcReadPort_0_1_prd = rat_5_prfIdx;
      5'b00110 : _zz_io_srcReadPort_0_1_prd = rat_6_prfIdx;
      5'b00111 : _zz_io_srcReadPort_0_1_prd = rat_7_prfIdx;
      5'b01000 : _zz_io_srcReadPort_0_1_prd = rat_8_prfIdx;
      5'b01001 : _zz_io_srcReadPort_0_1_prd = rat_9_prfIdx;
      5'b01010 : _zz_io_srcReadPort_0_1_prd = rat_10_prfIdx;
      5'b01011 : _zz_io_srcReadPort_0_1_prd = rat_11_prfIdx;
      5'b01100 : _zz_io_srcReadPort_0_1_prd = rat_12_prfIdx;
      5'b01101 : _zz_io_srcReadPort_0_1_prd = rat_13_prfIdx;
      5'b01110 : _zz_io_srcReadPort_0_1_prd = rat_14_prfIdx;
      5'b01111 : _zz_io_srcReadPort_0_1_prd = rat_15_prfIdx;
      5'b10000 : _zz_io_srcReadPort_0_1_prd = rat_16_prfIdx;
      5'b10001 : _zz_io_srcReadPort_0_1_prd = rat_17_prfIdx;
      5'b10010 : _zz_io_srcReadPort_0_1_prd = rat_18_prfIdx;
      5'b10011 : _zz_io_srcReadPort_0_1_prd = rat_19_prfIdx;
      5'b10100 : _zz_io_srcReadPort_0_1_prd = rat_20_prfIdx;
      5'b10101 : _zz_io_srcReadPort_0_1_prd = rat_21_prfIdx;
      5'b10110 : _zz_io_srcReadPort_0_1_prd = rat_22_prfIdx;
      5'b10111 : _zz_io_srcReadPort_0_1_prd = rat_23_prfIdx;
      5'b11000 : _zz_io_srcReadPort_0_1_prd = rat_24_prfIdx;
      5'b11001 : _zz_io_srcReadPort_0_1_prd = rat_25_prfIdx;
      5'b11010 : _zz_io_srcReadPort_0_1_prd = rat_26_prfIdx;
      5'b11011 : _zz_io_srcReadPort_0_1_prd = rat_27_prfIdx;
      5'b11100 : _zz_io_srcReadPort_0_1_prd = rat_28_prfIdx;
      5'b11101 : _zz_io_srcReadPort_0_1_prd = rat_29_prfIdx;
      5'b11110 : _zz_io_srcReadPort_0_1_prd = rat_30_prfIdx;
      default : _zz_io_srcReadPort_0_1_prd = rat_31_prfIdx;
    endcase
  end

  always @(*) begin
    case(_zz_io_srcReadPort_0_1_valid_1)
      5'b00000 : _zz_io_srcReadPort_0_1_valid = rat_0_valid;
      5'b00001 : _zz_io_srcReadPort_0_1_valid = rat_1_valid;
      5'b00010 : _zz_io_srcReadPort_0_1_valid = rat_2_valid;
      5'b00011 : _zz_io_srcReadPort_0_1_valid = rat_3_valid;
      5'b00100 : _zz_io_srcReadPort_0_1_valid = rat_4_valid;
      5'b00101 : _zz_io_srcReadPort_0_1_valid = rat_5_valid;
      5'b00110 : _zz_io_srcReadPort_0_1_valid = rat_6_valid;
      5'b00111 : _zz_io_srcReadPort_0_1_valid = rat_7_valid;
      5'b01000 : _zz_io_srcReadPort_0_1_valid = rat_8_valid;
      5'b01001 : _zz_io_srcReadPort_0_1_valid = rat_9_valid;
      5'b01010 : _zz_io_srcReadPort_0_1_valid = rat_10_valid;
      5'b01011 : _zz_io_srcReadPort_0_1_valid = rat_11_valid;
      5'b01100 : _zz_io_srcReadPort_0_1_valid = rat_12_valid;
      5'b01101 : _zz_io_srcReadPort_0_1_valid = rat_13_valid;
      5'b01110 : _zz_io_srcReadPort_0_1_valid = rat_14_valid;
      5'b01111 : _zz_io_srcReadPort_0_1_valid = rat_15_valid;
      5'b10000 : _zz_io_srcReadPort_0_1_valid = rat_16_valid;
      5'b10001 : _zz_io_srcReadPort_0_1_valid = rat_17_valid;
      5'b10010 : _zz_io_srcReadPort_0_1_valid = rat_18_valid;
      5'b10011 : _zz_io_srcReadPort_0_1_valid = rat_19_valid;
      5'b10100 : _zz_io_srcReadPort_0_1_valid = rat_20_valid;
      5'b10101 : _zz_io_srcReadPort_0_1_valid = rat_21_valid;
      5'b10110 : _zz_io_srcReadPort_0_1_valid = rat_22_valid;
      5'b10111 : _zz_io_srcReadPort_0_1_valid = rat_23_valid;
      5'b11000 : _zz_io_srcReadPort_0_1_valid = rat_24_valid;
      5'b11001 : _zz_io_srcReadPort_0_1_valid = rat_25_valid;
      5'b11010 : _zz_io_srcReadPort_0_1_valid = rat_26_valid;
      5'b11011 : _zz_io_srcReadPort_0_1_valid = rat_27_valid;
      5'b11100 : _zz_io_srcReadPort_0_1_valid = rat_28_valid;
      5'b11101 : _zz_io_srcReadPort_0_1_valid = rat_29_valid;
      5'b11110 : _zz_io_srcReadPort_0_1_valid = rat_30_valid;
      default : _zz_io_srcReadPort_0_1_valid = rat_31_valid;
    endcase
  end

  always @(*) begin
    case(_zz_io_srcReadPort_1_0_prd_1)
      5'b00000 : _zz_io_srcReadPort_1_0_prd = rat_0_prfIdx;
      5'b00001 : _zz_io_srcReadPort_1_0_prd = rat_1_prfIdx;
      5'b00010 : _zz_io_srcReadPort_1_0_prd = rat_2_prfIdx;
      5'b00011 : _zz_io_srcReadPort_1_0_prd = rat_3_prfIdx;
      5'b00100 : _zz_io_srcReadPort_1_0_prd = rat_4_prfIdx;
      5'b00101 : _zz_io_srcReadPort_1_0_prd = rat_5_prfIdx;
      5'b00110 : _zz_io_srcReadPort_1_0_prd = rat_6_prfIdx;
      5'b00111 : _zz_io_srcReadPort_1_0_prd = rat_7_prfIdx;
      5'b01000 : _zz_io_srcReadPort_1_0_prd = rat_8_prfIdx;
      5'b01001 : _zz_io_srcReadPort_1_0_prd = rat_9_prfIdx;
      5'b01010 : _zz_io_srcReadPort_1_0_prd = rat_10_prfIdx;
      5'b01011 : _zz_io_srcReadPort_1_0_prd = rat_11_prfIdx;
      5'b01100 : _zz_io_srcReadPort_1_0_prd = rat_12_prfIdx;
      5'b01101 : _zz_io_srcReadPort_1_0_prd = rat_13_prfIdx;
      5'b01110 : _zz_io_srcReadPort_1_0_prd = rat_14_prfIdx;
      5'b01111 : _zz_io_srcReadPort_1_0_prd = rat_15_prfIdx;
      5'b10000 : _zz_io_srcReadPort_1_0_prd = rat_16_prfIdx;
      5'b10001 : _zz_io_srcReadPort_1_0_prd = rat_17_prfIdx;
      5'b10010 : _zz_io_srcReadPort_1_0_prd = rat_18_prfIdx;
      5'b10011 : _zz_io_srcReadPort_1_0_prd = rat_19_prfIdx;
      5'b10100 : _zz_io_srcReadPort_1_0_prd = rat_20_prfIdx;
      5'b10101 : _zz_io_srcReadPort_1_0_prd = rat_21_prfIdx;
      5'b10110 : _zz_io_srcReadPort_1_0_prd = rat_22_prfIdx;
      5'b10111 : _zz_io_srcReadPort_1_0_prd = rat_23_prfIdx;
      5'b11000 : _zz_io_srcReadPort_1_0_prd = rat_24_prfIdx;
      5'b11001 : _zz_io_srcReadPort_1_0_prd = rat_25_prfIdx;
      5'b11010 : _zz_io_srcReadPort_1_0_prd = rat_26_prfIdx;
      5'b11011 : _zz_io_srcReadPort_1_0_prd = rat_27_prfIdx;
      5'b11100 : _zz_io_srcReadPort_1_0_prd = rat_28_prfIdx;
      5'b11101 : _zz_io_srcReadPort_1_0_prd = rat_29_prfIdx;
      5'b11110 : _zz_io_srcReadPort_1_0_prd = rat_30_prfIdx;
      default : _zz_io_srcReadPort_1_0_prd = rat_31_prfIdx;
    endcase
  end

  always @(*) begin
    case(_zz_io_srcReadPort_1_0_valid_1)
      5'b00000 : _zz_io_srcReadPort_1_0_valid = rat_0_valid;
      5'b00001 : _zz_io_srcReadPort_1_0_valid = rat_1_valid;
      5'b00010 : _zz_io_srcReadPort_1_0_valid = rat_2_valid;
      5'b00011 : _zz_io_srcReadPort_1_0_valid = rat_3_valid;
      5'b00100 : _zz_io_srcReadPort_1_0_valid = rat_4_valid;
      5'b00101 : _zz_io_srcReadPort_1_0_valid = rat_5_valid;
      5'b00110 : _zz_io_srcReadPort_1_0_valid = rat_6_valid;
      5'b00111 : _zz_io_srcReadPort_1_0_valid = rat_7_valid;
      5'b01000 : _zz_io_srcReadPort_1_0_valid = rat_8_valid;
      5'b01001 : _zz_io_srcReadPort_1_0_valid = rat_9_valid;
      5'b01010 : _zz_io_srcReadPort_1_0_valid = rat_10_valid;
      5'b01011 : _zz_io_srcReadPort_1_0_valid = rat_11_valid;
      5'b01100 : _zz_io_srcReadPort_1_0_valid = rat_12_valid;
      5'b01101 : _zz_io_srcReadPort_1_0_valid = rat_13_valid;
      5'b01110 : _zz_io_srcReadPort_1_0_valid = rat_14_valid;
      5'b01111 : _zz_io_srcReadPort_1_0_valid = rat_15_valid;
      5'b10000 : _zz_io_srcReadPort_1_0_valid = rat_16_valid;
      5'b10001 : _zz_io_srcReadPort_1_0_valid = rat_17_valid;
      5'b10010 : _zz_io_srcReadPort_1_0_valid = rat_18_valid;
      5'b10011 : _zz_io_srcReadPort_1_0_valid = rat_19_valid;
      5'b10100 : _zz_io_srcReadPort_1_0_valid = rat_20_valid;
      5'b10101 : _zz_io_srcReadPort_1_0_valid = rat_21_valid;
      5'b10110 : _zz_io_srcReadPort_1_0_valid = rat_22_valid;
      5'b10111 : _zz_io_srcReadPort_1_0_valid = rat_23_valid;
      5'b11000 : _zz_io_srcReadPort_1_0_valid = rat_24_valid;
      5'b11001 : _zz_io_srcReadPort_1_0_valid = rat_25_valid;
      5'b11010 : _zz_io_srcReadPort_1_0_valid = rat_26_valid;
      5'b11011 : _zz_io_srcReadPort_1_0_valid = rat_27_valid;
      5'b11100 : _zz_io_srcReadPort_1_0_valid = rat_28_valid;
      5'b11101 : _zz_io_srcReadPort_1_0_valid = rat_29_valid;
      5'b11110 : _zz_io_srcReadPort_1_0_valid = rat_30_valid;
      default : _zz_io_srcReadPort_1_0_valid = rat_31_valid;
    endcase
  end

  always @(*) begin
    case(_zz_io_srcReadPort_1_1_prd_1)
      5'b00000 : _zz_io_srcReadPort_1_1_prd = rat_0_prfIdx;
      5'b00001 : _zz_io_srcReadPort_1_1_prd = rat_1_prfIdx;
      5'b00010 : _zz_io_srcReadPort_1_1_prd = rat_2_prfIdx;
      5'b00011 : _zz_io_srcReadPort_1_1_prd = rat_3_prfIdx;
      5'b00100 : _zz_io_srcReadPort_1_1_prd = rat_4_prfIdx;
      5'b00101 : _zz_io_srcReadPort_1_1_prd = rat_5_prfIdx;
      5'b00110 : _zz_io_srcReadPort_1_1_prd = rat_6_prfIdx;
      5'b00111 : _zz_io_srcReadPort_1_1_prd = rat_7_prfIdx;
      5'b01000 : _zz_io_srcReadPort_1_1_prd = rat_8_prfIdx;
      5'b01001 : _zz_io_srcReadPort_1_1_prd = rat_9_prfIdx;
      5'b01010 : _zz_io_srcReadPort_1_1_prd = rat_10_prfIdx;
      5'b01011 : _zz_io_srcReadPort_1_1_prd = rat_11_prfIdx;
      5'b01100 : _zz_io_srcReadPort_1_1_prd = rat_12_prfIdx;
      5'b01101 : _zz_io_srcReadPort_1_1_prd = rat_13_prfIdx;
      5'b01110 : _zz_io_srcReadPort_1_1_prd = rat_14_prfIdx;
      5'b01111 : _zz_io_srcReadPort_1_1_prd = rat_15_prfIdx;
      5'b10000 : _zz_io_srcReadPort_1_1_prd = rat_16_prfIdx;
      5'b10001 : _zz_io_srcReadPort_1_1_prd = rat_17_prfIdx;
      5'b10010 : _zz_io_srcReadPort_1_1_prd = rat_18_prfIdx;
      5'b10011 : _zz_io_srcReadPort_1_1_prd = rat_19_prfIdx;
      5'b10100 : _zz_io_srcReadPort_1_1_prd = rat_20_prfIdx;
      5'b10101 : _zz_io_srcReadPort_1_1_prd = rat_21_prfIdx;
      5'b10110 : _zz_io_srcReadPort_1_1_prd = rat_22_prfIdx;
      5'b10111 : _zz_io_srcReadPort_1_1_prd = rat_23_prfIdx;
      5'b11000 : _zz_io_srcReadPort_1_1_prd = rat_24_prfIdx;
      5'b11001 : _zz_io_srcReadPort_1_1_prd = rat_25_prfIdx;
      5'b11010 : _zz_io_srcReadPort_1_1_prd = rat_26_prfIdx;
      5'b11011 : _zz_io_srcReadPort_1_1_prd = rat_27_prfIdx;
      5'b11100 : _zz_io_srcReadPort_1_1_prd = rat_28_prfIdx;
      5'b11101 : _zz_io_srcReadPort_1_1_prd = rat_29_prfIdx;
      5'b11110 : _zz_io_srcReadPort_1_1_prd = rat_30_prfIdx;
      default : _zz_io_srcReadPort_1_1_prd = rat_31_prfIdx;
    endcase
  end

  always @(*) begin
    case(_zz_io_srcReadPort_1_1_valid_1)
      5'b00000 : _zz_io_srcReadPort_1_1_valid = rat_0_valid;
      5'b00001 : _zz_io_srcReadPort_1_1_valid = rat_1_valid;
      5'b00010 : _zz_io_srcReadPort_1_1_valid = rat_2_valid;
      5'b00011 : _zz_io_srcReadPort_1_1_valid = rat_3_valid;
      5'b00100 : _zz_io_srcReadPort_1_1_valid = rat_4_valid;
      5'b00101 : _zz_io_srcReadPort_1_1_valid = rat_5_valid;
      5'b00110 : _zz_io_srcReadPort_1_1_valid = rat_6_valid;
      5'b00111 : _zz_io_srcReadPort_1_1_valid = rat_7_valid;
      5'b01000 : _zz_io_srcReadPort_1_1_valid = rat_8_valid;
      5'b01001 : _zz_io_srcReadPort_1_1_valid = rat_9_valid;
      5'b01010 : _zz_io_srcReadPort_1_1_valid = rat_10_valid;
      5'b01011 : _zz_io_srcReadPort_1_1_valid = rat_11_valid;
      5'b01100 : _zz_io_srcReadPort_1_1_valid = rat_12_valid;
      5'b01101 : _zz_io_srcReadPort_1_1_valid = rat_13_valid;
      5'b01110 : _zz_io_srcReadPort_1_1_valid = rat_14_valid;
      5'b01111 : _zz_io_srcReadPort_1_1_valid = rat_15_valid;
      5'b10000 : _zz_io_srcReadPort_1_1_valid = rat_16_valid;
      5'b10001 : _zz_io_srcReadPort_1_1_valid = rat_17_valid;
      5'b10010 : _zz_io_srcReadPort_1_1_valid = rat_18_valid;
      5'b10011 : _zz_io_srcReadPort_1_1_valid = rat_19_valid;
      5'b10100 : _zz_io_srcReadPort_1_1_valid = rat_20_valid;
      5'b10101 : _zz_io_srcReadPort_1_1_valid = rat_21_valid;
      5'b10110 : _zz_io_srcReadPort_1_1_valid = rat_22_valid;
      5'b10111 : _zz_io_srcReadPort_1_1_valid = rat_23_valid;
      5'b11000 : _zz_io_srcReadPort_1_1_valid = rat_24_valid;
      5'b11001 : _zz_io_srcReadPort_1_1_valid = rat_25_valid;
      5'b11010 : _zz_io_srcReadPort_1_1_valid = rat_26_valid;
      5'b11011 : _zz_io_srcReadPort_1_1_valid = rat_27_valid;
      5'b11100 : _zz_io_srcReadPort_1_1_valid = rat_28_valid;
      5'b11101 : _zz_io_srcReadPort_1_1_valid = rat_29_valid;
      5'b11110 : _zz_io_srcReadPort_1_1_valid = rat_30_valid;
      default : _zz_io_srcReadPort_1_1_valid = rat_31_valid;
    endcase
  end

  always @(*) begin
    case(_zz_io_prevPRDReadPort_0_prd_1)
      5'b00000 : _zz_io_prevPRDReadPort_0_prd = rat_0_prfIdx;
      5'b00001 : _zz_io_prevPRDReadPort_0_prd = rat_1_prfIdx;
      5'b00010 : _zz_io_prevPRDReadPort_0_prd = rat_2_prfIdx;
      5'b00011 : _zz_io_prevPRDReadPort_0_prd = rat_3_prfIdx;
      5'b00100 : _zz_io_prevPRDReadPort_0_prd = rat_4_prfIdx;
      5'b00101 : _zz_io_prevPRDReadPort_0_prd = rat_5_prfIdx;
      5'b00110 : _zz_io_prevPRDReadPort_0_prd = rat_6_prfIdx;
      5'b00111 : _zz_io_prevPRDReadPort_0_prd = rat_7_prfIdx;
      5'b01000 : _zz_io_prevPRDReadPort_0_prd = rat_8_prfIdx;
      5'b01001 : _zz_io_prevPRDReadPort_0_prd = rat_9_prfIdx;
      5'b01010 : _zz_io_prevPRDReadPort_0_prd = rat_10_prfIdx;
      5'b01011 : _zz_io_prevPRDReadPort_0_prd = rat_11_prfIdx;
      5'b01100 : _zz_io_prevPRDReadPort_0_prd = rat_12_prfIdx;
      5'b01101 : _zz_io_prevPRDReadPort_0_prd = rat_13_prfIdx;
      5'b01110 : _zz_io_prevPRDReadPort_0_prd = rat_14_prfIdx;
      5'b01111 : _zz_io_prevPRDReadPort_0_prd = rat_15_prfIdx;
      5'b10000 : _zz_io_prevPRDReadPort_0_prd = rat_16_prfIdx;
      5'b10001 : _zz_io_prevPRDReadPort_0_prd = rat_17_prfIdx;
      5'b10010 : _zz_io_prevPRDReadPort_0_prd = rat_18_prfIdx;
      5'b10011 : _zz_io_prevPRDReadPort_0_prd = rat_19_prfIdx;
      5'b10100 : _zz_io_prevPRDReadPort_0_prd = rat_20_prfIdx;
      5'b10101 : _zz_io_prevPRDReadPort_0_prd = rat_21_prfIdx;
      5'b10110 : _zz_io_prevPRDReadPort_0_prd = rat_22_prfIdx;
      5'b10111 : _zz_io_prevPRDReadPort_0_prd = rat_23_prfIdx;
      5'b11000 : _zz_io_prevPRDReadPort_0_prd = rat_24_prfIdx;
      5'b11001 : _zz_io_prevPRDReadPort_0_prd = rat_25_prfIdx;
      5'b11010 : _zz_io_prevPRDReadPort_0_prd = rat_26_prfIdx;
      5'b11011 : _zz_io_prevPRDReadPort_0_prd = rat_27_prfIdx;
      5'b11100 : _zz_io_prevPRDReadPort_0_prd = rat_28_prfIdx;
      5'b11101 : _zz_io_prevPRDReadPort_0_prd = rat_29_prfIdx;
      5'b11110 : _zz_io_prevPRDReadPort_0_prd = rat_30_prfIdx;
      default : _zz_io_prevPRDReadPort_0_prd = rat_31_prfIdx;
    endcase
  end

  always @(*) begin
    case(_zz_io_prevPRDReadPort_0_valid_1)
      5'b00000 : _zz_io_prevPRDReadPort_0_valid = rat_0_valid;
      5'b00001 : _zz_io_prevPRDReadPort_0_valid = rat_1_valid;
      5'b00010 : _zz_io_prevPRDReadPort_0_valid = rat_2_valid;
      5'b00011 : _zz_io_prevPRDReadPort_0_valid = rat_3_valid;
      5'b00100 : _zz_io_prevPRDReadPort_0_valid = rat_4_valid;
      5'b00101 : _zz_io_prevPRDReadPort_0_valid = rat_5_valid;
      5'b00110 : _zz_io_prevPRDReadPort_0_valid = rat_6_valid;
      5'b00111 : _zz_io_prevPRDReadPort_0_valid = rat_7_valid;
      5'b01000 : _zz_io_prevPRDReadPort_0_valid = rat_8_valid;
      5'b01001 : _zz_io_prevPRDReadPort_0_valid = rat_9_valid;
      5'b01010 : _zz_io_prevPRDReadPort_0_valid = rat_10_valid;
      5'b01011 : _zz_io_prevPRDReadPort_0_valid = rat_11_valid;
      5'b01100 : _zz_io_prevPRDReadPort_0_valid = rat_12_valid;
      5'b01101 : _zz_io_prevPRDReadPort_0_valid = rat_13_valid;
      5'b01110 : _zz_io_prevPRDReadPort_0_valid = rat_14_valid;
      5'b01111 : _zz_io_prevPRDReadPort_0_valid = rat_15_valid;
      5'b10000 : _zz_io_prevPRDReadPort_0_valid = rat_16_valid;
      5'b10001 : _zz_io_prevPRDReadPort_0_valid = rat_17_valid;
      5'b10010 : _zz_io_prevPRDReadPort_0_valid = rat_18_valid;
      5'b10011 : _zz_io_prevPRDReadPort_0_valid = rat_19_valid;
      5'b10100 : _zz_io_prevPRDReadPort_0_valid = rat_20_valid;
      5'b10101 : _zz_io_prevPRDReadPort_0_valid = rat_21_valid;
      5'b10110 : _zz_io_prevPRDReadPort_0_valid = rat_22_valid;
      5'b10111 : _zz_io_prevPRDReadPort_0_valid = rat_23_valid;
      5'b11000 : _zz_io_prevPRDReadPort_0_valid = rat_24_valid;
      5'b11001 : _zz_io_prevPRDReadPort_0_valid = rat_25_valid;
      5'b11010 : _zz_io_prevPRDReadPort_0_valid = rat_26_valid;
      5'b11011 : _zz_io_prevPRDReadPort_0_valid = rat_27_valid;
      5'b11100 : _zz_io_prevPRDReadPort_0_valid = rat_28_valid;
      5'b11101 : _zz_io_prevPRDReadPort_0_valid = rat_29_valid;
      5'b11110 : _zz_io_prevPRDReadPort_0_valid = rat_30_valid;
      default : _zz_io_prevPRDReadPort_0_valid = rat_31_valid;
    endcase
  end

  always @(*) begin
    case(_zz_io_prevPRDReadPort_1_prd_1)
      5'b00000 : _zz_io_prevPRDReadPort_1_prd = rat_0_prfIdx;
      5'b00001 : _zz_io_prevPRDReadPort_1_prd = rat_1_prfIdx;
      5'b00010 : _zz_io_prevPRDReadPort_1_prd = rat_2_prfIdx;
      5'b00011 : _zz_io_prevPRDReadPort_1_prd = rat_3_prfIdx;
      5'b00100 : _zz_io_prevPRDReadPort_1_prd = rat_4_prfIdx;
      5'b00101 : _zz_io_prevPRDReadPort_1_prd = rat_5_prfIdx;
      5'b00110 : _zz_io_prevPRDReadPort_1_prd = rat_6_prfIdx;
      5'b00111 : _zz_io_prevPRDReadPort_1_prd = rat_7_prfIdx;
      5'b01000 : _zz_io_prevPRDReadPort_1_prd = rat_8_prfIdx;
      5'b01001 : _zz_io_prevPRDReadPort_1_prd = rat_9_prfIdx;
      5'b01010 : _zz_io_prevPRDReadPort_1_prd = rat_10_prfIdx;
      5'b01011 : _zz_io_prevPRDReadPort_1_prd = rat_11_prfIdx;
      5'b01100 : _zz_io_prevPRDReadPort_1_prd = rat_12_prfIdx;
      5'b01101 : _zz_io_prevPRDReadPort_1_prd = rat_13_prfIdx;
      5'b01110 : _zz_io_prevPRDReadPort_1_prd = rat_14_prfIdx;
      5'b01111 : _zz_io_prevPRDReadPort_1_prd = rat_15_prfIdx;
      5'b10000 : _zz_io_prevPRDReadPort_1_prd = rat_16_prfIdx;
      5'b10001 : _zz_io_prevPRDReadPort_1_prd = rat_17_prfIdx;
      5'b10010 : _zz_io_prevPRDReadPort_1_prd = rat_18_prfIdx;
      5'b10011 : _zz_io_prevPRDReadPort_1_prd = rat_19_prfIdx;
      5'b10100 : _zz_io_prevPRDReadPort_1_prd = rat_20_prfIdx;
      5'b10101 : _zz_io_prevPRDReadPort_1_prd = rat_21_prfIdx;
      5'b10110 : _zz_io_prevPRDReadPort_1_prd = rat_22_prfIdx;
      5'b10111 : _zz_io_prevPRDReadPort_1_prd = rat_23_prfIdx;
      5'b11000 : _zz_io_prevPRDReadPort_1_prd = rat_24_prfIdx;
      5'b11001 : _zz_io_prevPRDReadPort_1_prd = rat_25_prfIdx;
      5'b11010 : _zz_io_prevPRDReadPort_1_prd = rat_26_prfIdx;
      5'b11011 : _zz_io_prevPRDReadPort_1_prd = rat_27_prfIdx;
      5'b11100 : _zz_io_prevPRDReadPort_1_prd = rat_28_prfIdx;
      5'b11101 : _zz_io_prevPRDReadPort_1_prd = rat_29_prfIdx;
      5'b11110 : _zz_io_prevPRDReadPort_1_prd = rat_30_prfIdx;
      default : _zz_io_prevPRDReadPort_1_prd = rat_31_prfIdx;
    endcase
  end

  always @(*) begin
    case(_zz_io_prevPRDReadPort_1_valid_1)
      5'b00000 : _zz_io_prevPRDReadPort_1_valid = rat_0_valid;
      5'b00001 : _zz_io_prevPRDReadPort_1_valid = rat_1_valid;
      5'b00010 : _zz_io_prevPRDReadPort_1_valid = rat_2_valid;
      5'b00011 : _zz_io_prevPRDReadPort_1_valid = rat_3_valid;
      5'b00100 : _zz_io_prevPRDReadPort_1_valid = rat_4_valid;
      5'b00101 : _zz_io_prevPRDReadPort_1_valid = rat_5_valid;
      5'b00110 : _zz_io_prevPRDReadPort_1_valid = rat_6_valid;
      5'b00111 : _zz_io_prevPRDReadPort_1_valid = rat_7_valid;
      5'b01000 : _zz_io_prevPRDReadPort_1_valid = rat_8_valid;
      5'b01001 : _zz_io_prevPRDReadPort_1_valid = rat_9_valid;
      5'b01010 : _zz_io_prevPRDReadPort_1_valid = rat_10_valid;
      5'b01011 : _zz_io_prevPRDReadPort_1_valid = rat_11_valid;
      5'b01100 : _zz_io_prevPRDReadPort_1_valid = rat_12_valid;
      5'b01101 : _zz_io_prevPRDReadPort_1_valid = rat_13_valid;
      5'b01110 : _zz_io_prevPRDReadPort_1_valid = rat_14_valid;
      5'b01111 : _zz_io_prevPRDReadPort_1_valid = rat_15_valid;
      5'b10000 : _zz_io_prevPRDReadPort_1_valid = rat_16_valid;
      5'b10001 : _zz_io_prevPRDReadPort_1_valid = rat_17_valid;
      5'b10010 : _zz_io_prevPRDReadPort_1_valid = rat_18_valid;
      5'b10011 : _zz_io_prevPRDReadPort_1_valid = rat_19_valid;
      5'b10100 : _zz_io_prevPRDReadPort_1_valid = rat_20_valid;
      5'b10101 : _zz_io_prevPRDReadPort_1_valid = rat_21_valid;
      5'b10110 : _zz_io_prevPRDReadPort_1_valid = rat_22_valid;
      5'b10111 : _zz_io_prevPRDReadPort_1_valid = rat_23_valid;
      5'b11000 : _zz_io_prevPRDReadPort_1_valid = rat_24_valid;
      5'b11001 : _zz_io_prevPRDReadPort_1_valid = rat_25_valid;
      5'b11010 : _zz_io_prevPRDReadPort_1_valid = rat_26_valid;
      5'b11011 : _zz_io_prevPRDReadPort_1_valid = rat_27_valid;
      5'b11100 : _zz_io_prevPRDReadPort_1_valid = rat_28_valid;
      5'b11101 : _zz_io_prevPRDReadPort_1_valid = rat_29_valid;
      5'b11110 : _zz_io_prevPRDReadPort_1_valid = rat_30_valid;
      default : _zz_io_prevPRDReadPort_1_valid = rat_31_valid;
    endcase
  end

  assign when_RAT_l30 = (io_updatePort_0_wen && (rat_0_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_1 = (io_updatePort_1_wen && (rat_0_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_2 = (io_updatePort_2_wen && (rat_0_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_3 = (io_updatePort_3_wen && (rat_0_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_4 = (io_updatePort_4_wen && (rat_0_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_5 = (io_updatePort_0_wen && (rat_1_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_6 = (io_updatePort_1_wen && (rat_1_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_7 = (io_updatePort_2_wen && (rat_1_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_8 = (io_updatePort_3_wen && (rat_1_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_9 = (io_updatePort_4_wen && (rat_1_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_10 = (io_updatePort_0_wen && (rat_2_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_11 = (io_updatePort_1_wen && (rat_2_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_12 = (io_updatePort_2_wen && (rat_2_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_13 = (io_updatePort_3_wen && (rat_2_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_14 = (io_updatePort_4_wen && (rat_2_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_15 = (io_updatePort_0_wen && (rat_3_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_16 = (io_updatePort_1_wen && (rat_3_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_17 = (io_updatePort_2_wen && (rat_3_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_18 = (io_updatePort_3_wen && (rat_3_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_19 = (io_updatePort_4_wen && (rat_3_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_20 = (io_updatePort_0_wen && (rat_4_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_21 = (io_updatePort_1_wen && (rat_4_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_22 = (io_updatePort_2_wen && (rat_4_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_23 = (io_updatePort_3_wen && (rat_4_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_24 = (io_updatePort_4_wen && (rat_4_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_25 = (io_updatePort_0_wen && (rat_5_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_26 = (io_updatePort_1_wen && (rat_5_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_27 = (io_updatePort_2_wen && (rat_5_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_28 = (io_updatePort_3_wen && (rat_5_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_29 = (io_updatePort_4_wen && (rat_5_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_30 = (io_updatePort_0_wen && (rat_6_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_31 = (io_updatePort_1_wen && (rat_6_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_32 = (io_updatePort_2_wen && (rat_6_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_33 = (io_updatePort_3_wen && (rat_6_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_34 = (io_updatePort_4_wen && (rat_6_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_35 = (io_updatePort_0_wen && (rat_7_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_36 = (io_updatePort_1_wen && (rat_7_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_37 = (io_updatePort_2_wen && (rat_7_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_38 = (io_updatePort_3_wen && (rat_7_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_39 = (io_updatePort_4_wen && (rat_7_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_40 = (io_updatePort_0_wen && (rat_8_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_41 = (io_updatePort_1_wen && (rat_8_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_42 = (io_updatePort_2_wen && (rat_8_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_43 = (io_updatePort_3_wen && (rat_8_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_44 = (io_updatePort_4_wen && (rat_8_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_45 = (io_updatePort_0_wen && (rat_9_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_46 = (io_updatePort_1_wen && (rat_9_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_47 = (io_updatePort_2_wen && (rat_9_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_48 = (io_updatePort_3_wen && (rat_9_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_49 = (io_updatePort_4_wen && (rat_9_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_50 = (io_updatePort_0_wen && (rat_10_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_51 = (io_updatePort_1_wen && (rat_10_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_52 = (io_updatePort_2_wen && (rat_10_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_53 = (io_updatePort_3_wen && (rat_10_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_54 = (io_updatePort_4_wen && (rat_10_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_55 = (io_updatePort_0_wen && (rat_11_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_56 = (io_updatePort_1_wen && (rat_11_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_57 = (io_updatePort_2_wen && (rat_11_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_58 = (io_updatePort_3_wen && (rat_11_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_59 = (io_updatePort_4_wen && (rat_11_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_60 = (io_updatePort_0_wen && (rat_12_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_61 = (io_updatePort_1_wen && (rat_12_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_62 = (io_updatePort_2_wen && (rat_12_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_63 = (io_updatePort_3_wen && (rat_12_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_64 = (io_updatePort_4_wen && (rat_12_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_65 = (io_updatePort_0_wen && (rat_13_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_66 = (io_updatePort_1_wen && (rat_13_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_67 = (io_updatePort_2_wen && (rat_13_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_68 = (io_updatePort_3_wen && (rat_13_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_69 = (io_updatePort_4_wen && (rat_13_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_70 = (io_updatePort_0_wen && (rat_14_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_71 = (io_updatePort_1_wen && (rat_14_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_72 = (io_updatePort_2_wen && (rat_14_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_73 = (io_updatePort_3_wen && (rat_14_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_74 = (io_updatePort_4_wen && (rat_14_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_75 = (io_updatePort_0_wen && (rat_15_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_76 = (io_updatePort_1_wen && (rat_15_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_77 = (io_updatePort_2_wen && (rat_15_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_78 = (io_updatePort_3_wen && (rat_15_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_79 = (io_updatePort_4_wen && (rat_15_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_80 = (io_updatePort_0_wen && (rat_16_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_81 = (io_updatePort_1_wen && (rat_16_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_82 = (io_updatePort_2_wen && (rat_16_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_83 = (io_updatePort_3_wen && (rat_16_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_84 = (io_updatePort_4_wen && (rat_16_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_85 = (io_updatePort_0_wen && (rat_17_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_86 = (io_updatePort_1_wen && (rat_17_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_87 = (io_updatePort_2_wen && (rat_17_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_88 = (io_updatePort_3_wen && (rat_17_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_89 = (io_updatePort_4_wen && (rat_17_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_90 = (io_updatePort_0_wen && (rat_18_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_91 = (io_updatePort_1_wen && (rat_18_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_92 = (io_updatePort_2_wen && (rat_18_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_93 = (io_updatePort_3_wen && (rat_18_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_94 = (io_updatePort_4_wen && (rat_18_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_95 = (io_updatePort_0_wen && (rat_19_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_96 = (io_updatePort_1_wen && (rat_19_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_97 = (io_updatePort_2_wen && (rat_19_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_98 = (io_updatePort_3_wen && (rat_19_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_99 = (io_updatePort_4_wen && (rat_19_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_100 = (io_updatePort_0_wen && (rat_20_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_101 = (io_updatePort_1_wen && (rat_20_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_102 = (io_updatePort_2_wen && (rat_20_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_103 = (io_updatePort_3_wen && (rat_20_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_104 = (io_updatePort_4_wen && (rat_20_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_105 = (io_updatePort_0_wen && (rat_21_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_106 = (io_updatePort_1_wen && (rat_21_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_107 = (io_updatePort_2_wen && (rat_21_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_108 = (io_updatePort_3_wen && (rat_21_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_109 = (io_updatePort_4_wen && (rat_21_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_110 = (io_updatePort_0_wen && (rat_22_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_111 = (io_updatePort_1_wen && (rat_22_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_112 = (io_updatePort_2_wen && (rat_22_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_113 = (io_updatePort_3_wen && (rat_22_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_114 = (io_updatePort_4_wen && (rat_22_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_115 = (io_updatePort_0_wen && (rat_23_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_116 = (io_updatePort_1_wen && (rat_23_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_117 = (io_updatePort_2_wen && (rat_23_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_118 = (io_updatePort_3_wen && (rat_23_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_119 = (io_updatePort_4_wen && (rat_23_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_120 = (io_updatePort_0_wen && (rat_24_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_121 = (io_updatePort_1_wen && (rat_24_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_122 = (io_updatePort_2_wen && (rat_24_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_123 = (io_updatePort_3_wen && (rat_24_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_124 = (io_updatePort_4_wen && (rat_24_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_125 = (io_updatePort_0_wen && (rat_25_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_126 = (io_updatePort_1_wen && (rat_25_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_127 = (io_updatePort_2_wen && (rat_25_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_128 = (io_updatePort_3_wen && (rat_25_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_129 = (io_updatePort_4_wen && (rat_25_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_130 = (io_updatePort_0_wen && (rat_26_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_131 = (io_updatePort_1_wen && (rat_26_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_132 = (io_updatePort_2_wen && (rat_26_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_133 = (io_updatePort_3_wen && (rat_26_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_134 = (io_updatePort_4_wen && (rat_26_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_135 = (io_updatePort_0_wen && (rat_27_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_136 = (io_updatePort_1_wen && (rat_27_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_137 = (io_updatePort_2_wen && (rat_27_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_138 = (io_updatePort_3_wen && (rat_27_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_139 = (io_updatePort_4_wen && (rat_27_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_140 = (io_updatePort_0_wen && (rat_28_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_141 = (io_updatePort_1_wen && (rat_28_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_142 = (io_updatePort_2_wen && (rat_28_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_143 = (io_updatePort_3_wen && (rat_28_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_144 = (io_updatePort_4_wen && (rat_28_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_145 = (io_updatePort_0_wen && (rat_29_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_146 = (io_updatePort_1_wen && (rat_29_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_147 = (io_updatePort_2_wen && (rat_29_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_148 = (io_updatePort_3_wen && (rat_29_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_149 = (io_updatePort_4_wen && (rat_29_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_150 = (io_updatePort_0_wen && (rat_30_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_151 = (io_updatePort_1_wen && (rat_30_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_152 = (io_updatePort_2_wen && (rat_30_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_153 = (io_updatePort_3_wen && (rat_30_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_154 = (io_updatePort_4_wen && (rat_30_prfIdx == io_updatePort_4_prd));
  assign when_RAT_l30_155 = (io_updatePort_0_wen && (rat_31_prfIdx == io_updatePort_0_prd));
  assign when_RAT_l30_156 = (io_updatePort_1_wen && (rat_31_prfIdx == io_updatePort_1_prd));
  assign when_RAT_l30_157 = (io_updatePort_2_wen && (rat_31_prfIdx == io_updatePort_2_prd));
  assign when_RAT_l30_158 = (io_updatePort_3_wen && (rat_31_prfIdx == io_updatePort_3_prd));
  assign when_RAT_l30_159 = (io_updatePort_4_wen && (rat_31_prfIdx == io_updatePort_4_prd));
  assign _zz_1 = ({31'd0,1'b1} <<< io_writePort_0_ard);
  assign _zz_2 = ({31'd0,1'b1} <<< io_writePort_0_ard);
  assign _zz_3 = ({31'd0,1'b1} <<< io_writePort_1_ard);
  assign _zz_4 = ({31'd0,1'b1} <<< io_writePort_1_ard);
  assign io_srcReadPort_0_0_prd = _zz_io_srcReadPort_0_0_prd;
  assign io_srcReadPort_0_0_valid = _zz_io_srcReadPort_0_0_valid;
  assign io_srcReadPort_0_1_prd = _zz_io_srcReadPort_0_1_prd;
  assign io_srcReadPort_0_1_valid = _zz_io_srcReadPort_0_1_valid;
  assign io_srcReadPort_1_0_prd = _zz_io_srcReadPort_1_0_prd;
  assign io_srcReadPort_1_0_valid = _zz_io_srcReadPort_1_0_valid;
  assign io_srcReadPort_1_1_prd = _zz_io_srcReadPort_1_1_prd;
  assign io_srcReadPort_1_1_valid = _zz_io_srcReadPort_1_1_valid;
  assign io_prevPRDReadPort_0_prd = _zz_io_prevPRDReadPort_0_prd;
  assign io_prevPRDReadPort_0_valid = _zz_io_prevPRDReadPort_0_valid;
  assign io_prevPRDReadPort_1_prd = _zz_io_prevPRDReadPort_1_prd;
  assign io_prevPRDReadPort_1_valid = _zz_io_prevPRDReadPort_1_valid;
  always @(posedge aclk) begin
    if(!aresetn) begin
      rat_0_prfIdx <= {5'd0, _zz_rat_0_prfIdx};
      rat_0_valid <= 1'b1;
      rat_1_prfIdx <= {5'd0, _zz_rat_1_prfIdx};
      rat_1_valid <= 1'b1;
      rat_2_prfIdx <= {5'd0, _zz_rat_2_prfIdx};
      rat_2_valid <= 1'b1;
      rat_3_prfIdx <= {5'd0, _zz_rat_3_prfIdx};
      rat_3_valid <= 1'b1;
      rat_4_prfIdx <= {5'd0, _zz_rat_4_prfIdx};
      rat_4_valid <= 1'b1;
      rat_5_prfIdx <= {5'd0, _zz_rat_5_prfIdx};
      rat_5_valid <= 1'b1;
      rat_6_prfIdx <= {5'd0, _zz_rat_6_prfIdx};
      rat_6_valid <= 1'b1;
      rat_7_prfIdx <= {5'd0, _zz_rat_7_prfIdx};
      rat_7_valid <= 1'b1;
      rat_8_prfIdx <= {5'd0, _zz_rat_8_prfIdx};
      rat_8_valid <= 1'b1;
      rat_9_prfIdx <= {5'd0, _zz_rat_9_prfIdx};
      rat_9_valid <= 1'b1;
      rat_10_prfIdx <= {5'd0, _zz_rat_10_prfIdx};
      rat_10_valid <= 1'b1;
      rat_11_prfIdx <= {5'd0, _zz_rat_11_prfIdx};
      rat_11_valid <= 1'b1;
      rat_12_prfIdx <= {5'd0, _zz_rat_12_prfIdx};
      rat_12_valid <= 1'b1;
      rat_13_prfIdx <= {5'd0, _zz_rat_13_prfIdx};
      rat_13_valid <= 1'b1;
      rat_14_prfIdx <= {5'd0, _zz_rat_14_prfIdx};
      rat_14_valid <= 1'b1;
      rat_15_prfIdx <= {5'd0, _zz_rat_15_prfIdx};
      rat_15_valid <= 1'b1;
      rat_16_prfIdx <= {5'd0, _zz_rat_16_prfIdx};
      rat_16_valid <= 1'b1;
      rat_17_prfIdx <= {5'd0, _zz_rat_17_prfIdx};
      rat_17_valid <= 1'b1;
      rat_18_prfIdx <= {5'd0, _zz_rat_18_prfIdx};
      rat_18_valid <= 1'b1;
      rat_19_prfIdx <= {5'd0, _zz_rat_19_prfIdx};
      rat_19_valid <= 1'b1;
      rat_20_prfIdx <= {5'd0, _zz_rat_20_prfIdx};
      rat_20_valid <= 1'b1;
      rat_21_prfIdx <= {5'd0, _zz_rat_21_prfIdx};
      rat_21_valid <= 1'b1;
      rat_22_prfIdx <= {5'd0, _zz_rat_22_prfIdx};
      rat_22_valid <= 1'b1;
      rat_23_prfIdx <= {5'd0, _zz_rat_23_prfIdx};
      rat_23_valid <= 1'b1;
      rat_24_prfIdx <= {5'd0, _zz_rat_24_prfIdx};
      rat_24_valid <= 1'b1;
      rat_25_prfIdx <= {5'd0, _zz_rat_25_prfIdx};
      rat_25_valid <= 1'b1;
      rat_26_prfIdx <= {5'd0, _zz_rat_26_prfIdx};
      rat_26_valid <= 1'b1;
      rat_27_prfIdx <= {5'd0, _zz_rat_27_prfIdx};
      rat_27_valid <= 1'b1;
      rat_28_prfIdx <= {5'd0, _zz_rat_28_prfIdx};
      rat_28_valid <= 1'b1;
      rat_29_prfIdx <= {5'd0, _zz_rat_29_prfIdx};
      rat_29_valid <= 1'b1;
      rat_30_prfIdx <= {5'd0, _zz_rat_30_prfIdx};
      rat_30_valid <= 1'b1;
      rat_31_prfIdx <= {5'd0, _zz_rat_31_prfIdx};
      rat_31_valid <= 1'b1;
    end else begin
      if(io_delayedRecovery) begin
        rat_0_prfIdx <= io_recoveryPort_0;
        rat_0_valid <= 1'b1;
        rat_1_prfIdx <= io_recoveryPort_1;
        rat_1_valid <= 1'b1;
        rat_2_prfIdx <= io_recoveryPort_2;
        rat_2_valid <= 1'b1;
        rat_3_prfIdx <= io_recoveryPort_3;
        rat_3_valid <= 1'b1;
        rat_4_prfIdx <= io_recoveryPort_4;
        rat_4_valid <= 1'b1;
        rat_5_prfIdx <= io_recoveryPort_5;
        rat_5_valid <= 1'b1;
        rat_6_prfIdx <= io_recoveryPort_6;
        rat_6_valid <= 1'b1;
        rat_7_prfIdx <= io_recoveryPort_7;
        rat_7_valid <= 1'b1;
        rat_8_prfIdx <= io_recoveryPort_8;
        rat_8_valid <= 1'b1;
        rat_9_prfIdx <= io_recoveryPort_9;
        rat_9_valid <= 1'b1;
        rat_10_prfIdx <= io_recoveryPort_10;
        rat_10_valid <= 1'b1;
        rat_11_prfIdx <= io_recoveryPort_11;
        rat_11_valid <= 1'b1;
        rat_12_prfIdx <= io_recoveryPort_12;
        rat_12_valid <= 1'b1;
        rat_13_prfIdx <= io_recoveryPort_13;
        rat_13_valid <= 1'b1;
        rat_14_prfIdx <= io_recoveryPort_14;
        rat_14_valid <= 1'b1;
        rat_15_prfIdx <= io_recoveryPort_15;
        rat_15_valid <= 1'b1;
        rat_16_prfIdx <= io_recoveryPort_16;
        rat_16_valid <= 1'b1;
        rat_17_prfIdx <= io_recoveryPort_17;
        rat_17_valid <= 1'b1;
        rat_18_prfIdx <= io_recoveryPort_18;
        rat_18_valid <= 1'b1;
        rat_19_prfIdx <= io_recoveryPort_19;
        rat_19_valid <= 1'b1;
        rat_20_prfIdx <= io_recoveryPort_20;
        rat_20_valid <= 1'b1;
        rat_21_prfIdx <= io_recoveryPort_21;
        rat_21_valid <= 1'b1;
        rat_22_prfIdx <= io_recoveryPort_22;
        rat_22_valid <= 1'b1;
        rat_23_prfIdx <= io_recoveryPort_23;
        rat_23_valid <= 1'b1;
        rat_24_prfIdx <= io_recoveryPort_24;
        rat_24_valid <= 1'b1;
        rat_25_prfIdx <= io_recoveryPort_25;
        rat_25_valid <= 1'b1;
        rat_26_prfIdx <= io_recoveryPort_26;
        rat_26_valid <= 1'b1;
        rat_27_prfIdx <= io_recoveryPort_27;
        rat_27_valid <= 1'b1;
        rat_28_prfIdx <= io_recoveryPort_28;
        rat_28_valid <= 1'b1;
        rat_29_prfIdx <= io_recoveryPort_29;
        rat_29_valid <= 1'b1;
        rat_30_prfIdx <= io_recoveryPort_30;
        rat_30_valid <= 1'b1;
        rat_31_prfIdx <= io_recoveryPort_31;
        rat_31_valid <= 1'b1;
      end else begin
        if(when_RAT_l30) begin
          rat_0_valid <= 1'b1;
        end
        if(when_RAT_l30_1) begin
          rat_0_valid <= 1'b1;
        end
        if(when_RAT_l30_2) begin
          rat_0_valid <= 1'b1;
        end
        if(when_RAT_l30_3) begin
          rat_0_valid <= 1'b1;
        end
        if(when_RAT_l30_4) begin
          rat_0_valid <= 1'b1;
        end
        if(when_RAT_l30_5) begin
          rat_1_valid <= 1'b1;
        end
        if(when_RAT_l30_6) begin
          rat_1_valid <= 1'b1;
        end
        if(when_RAT_l30_7) begin
          rat_1_valid <= 1'b1;
        end
        if(when_RAT_l30_8) begin
          rat_1_valid <= 1'b1;
        end
        if(when_RAT_l30_9) begin
          rat_1_valid <= 1'b1;
        end
        if(when_RAT_l30_10) begin
          rat_2_valid <= 1'b1;
        end
        if(when_RAT_l30_11) begin
          rat_2_valid <= 1'b1;
        end
        if(when_RAT_l30_12) begin
          rat_2_valid <= 1'b1;
        end
        if(when_RAT_l30_13) begin
          rat_2_valid <= 1'b1;
        end
        if(when_RAT_l30_14) begin
          rat_2_valid <= 1'b1;
        end
        if(when_RAT_l30_15) begin
          rat_3_valid <= 1'b1;
        end
        if(when_RAT_l30_16) begin
          rat_3_valid <= 1'b1;
        end
        if(when_RAT_l30_17) begin
          rat_3_valid <= 1'b1;
        end
        if(when_RAT_l30_18) begin
          rat_3_valid <= 1'b1;
        end
        if(when_RAT_l30_19) begin
          rat_3_valid <= 1'b1;
        end
        if(when_RAT_l30_20) begin
          rat_4_valid <= 1'b1;
        end
        if(when_RAT_l30_21) begin
          rat_4_valid <= 1'b1;
        end
        if(when_RAT_l30_22) begin
          rat_4_valid <= 1'b1;
        end
        if(when_RAT_l30_23) begin
          rat_4_valid <= 1'b1;
        end
        if(when_RAT_l30_24) begin
          rat_4_valid <= 1'b1;
        end
        if(when_RAT_l30_25) begin
          rat_5_valid <= 1'b1;
        end
        if(when_RAT_l30_26) begin
          rat_5_valid <= 1'b1;
        end
        if(when_RAT_l30_27) begin
          rat_5_valid <= 1'b1;
        end
        if(when_RAT_l30_28) begin
          rat_5_valid <= 1'b1;
        end
        if(when_RAT_l30_29) begin
          rat_5_valid <= 1'b1;
        end
        if(when_RAT_l30_30) begin
          rat_6_valid <= 1'b1;
        end
        if(when_RAT_l30_31) begin
          rat_6_valid <= 1'b1;
        end
        if(when_RAT_l30_32) begin
          rat_6_valid <= 1'b1;
        end
        if(when_RAT_l30_33) begin
          rat_6_valid <= 1'b1;
        end
        if(when_RAT_l30_34) begin
          rat_6_valid <= 1'b1;
        end
        if(when_RAT_l30_35) begin
          rat_7_valid <= 1'b1;
        end
        if(when_RAT_l30_36) begin
          rat_7_valid <= 1'b1;
        end
        if(when_RAT_l30_37) begin
          rat_7_valid <= 1'b1;
        end
        if(when_RAT_l30_38) begin
          rat_7_valid <= 1'b1;
        end
        if(when_RAT_l30_39) begin
          rat_7_valid <= 1'b1;
        end
        if(when_RAT_l30_40) begin
          rat_8_valid <= 1'b1;
        end
        if(when_RAT_l30_41) begin
          rat_8_valid <= 1'b1;
        end
        if(when_RAT_l30_42) begin
          rat_8_valid <= 1'b1;
        end
        if(when_RAT_l30_43) begin
          rat_8_valid <= 1'b1;
        end
        if(when_RAT_l30_44) begin
          rat_8_valid <= 1'b1;
        end
        if(when_RAT_l30_45) begin
          rat_9_valid <= 1'b1;
        end
        if(when_RAT_l30_46) begin
          rat_9_valid <= 1'b1;
        end
        if(when_RAT_l30_47) begin
          rat_9_valid <= 1'b1;
        end
        if(when_RAT_l30_48) begin
          rat_9_valid <= 1'b1;
        end
        if(when_RAT_l30_49) begin
          rat_9_valid <= 1'b1;
        end
        if(when_RAT_l30_50) begin
          rat_10_valid <= 1'b1;
        end
        if(when_RAT_l30_51) begin
          rat_10_valid <= 1'b1;
        end
        if(when_RAT_l30_52) begin
          rat_10_valid <= 1'b1;
        end
        if(when_RAT_l30_53) begin
          rat_10_valid <= 1'b1;
        end
        if(when_RAT_l30_54) begin
          rat_10_valid <= 1'b1;
        end
        if(when_RAT_l30_55) begin
          rat_11_valid <= 1'b1;
        end
        if(when_RAT_l30_56) begin
          rat_11_valid <= 1'b1;
        end
        if(when_RAT_l30_57) begin
          rat_11_valid <= 1'b1;
        end
        if(when_RAT_l30_58) begin
          rat_11_valid <= 1'b1;
        end
        if(when_RAT_l30_59) begin
          rat_11_valid <= 1'b1;
        end
        if(when_RAT_l30_60) begin
          rat_12_valid <= 1'b1;
        end
        if(when_RAT_l30_61) begin
          rat_12_valid <= 1'b1;
        end
        if(when_RAT_l30_62) begin
          rat_12_valid <= 1'b1;
        end
        if(when_RAT_l30_63) begin
          rat_12_valid <= 1'b1;
        end
        if(when_RAT_l30_64) begin
          rat_12_valid <= 1'b1;
        end
        if(when_RAT_l30_65) begin
          rat_13_valid <= 1'b1;
        end
        if(when_RAT_l30_66) begin
          rat_13_valid <= 1'b1;
        end
        if(when_RAT_l30_67) begin
          rat_13_valid <= 1'b1;
        end
        if(when_RAT_l30_68) begin
          rat_13_valid <= 1'b1;
        end
        if(when_RAT_l30_69) begin
          rat_13_valid <= 1'b1;
        end
        if(when_RAT_l30_70) begin
          rat_14_valid <= 1'b1;
        end
        if(when_RAT_l30_71) begin
          rat_14_valid <= 1'b1;
        end
        if(when_RAT_l30_72) begin
          rat_14_valid <= 1'b1;
        end
        if(when_RAT_l30_73) begin
          rat_14_valid <= 1'b1;
        end
        if(when_RAT_l30_74) begin
          rat_14_valid <= 1'b1;
        end
        if(when_RAT_l30_75) begin
          rat_15_valid <= 1'b1;
        end
        if(when_RAT_l30_76) begin
          rat_15_valid <= 1'b1;
        end
        if(when_RAT_l30_77) begin
          rat_15_valid <= 1'b1;
        end
        if(when_RAT_l30_78) begin
          rat_15_valid <= 1'b1;
        end
        if(when_RAT_l30_79) begin
          rat_15_valid <= 1'b1;
        end
        if(when_RAT_l30_80) begin
          rat_16_valid <= 1'b1;
        end
        if(when_RAT_l30_81) begin
          rat_16_valid <= 1'b1;
        end
        if(when_RAT_l30_82) begin
          rat_16_valid <= 1'b1;
        end
        if(when_RAT_l30_83) begin
          rat_16_valid <= 1'b1;
        end
        if(when_RAT_l30_84) begin
          rat_16_valid <= 1'b1;
        end
        if(when_RAT_l30_85) begin
          rat_17_valid <= 1'b1;
        end
        if(when_RAT_l30_86) begin
          rat_17_valid <= 1'b1;
        end
        if(when_RAT_l30_87) begin
          rat_17_valid <= 1'b1;
        end
        if(when_RAT_l30_88) begin
          rat_17_valid <= 1'b1;
        end
        if(when_RAT_l30_89) begin
          rat_17_valid <= 1'b1;
        end
        if(when_RAT_l30_90) begin
          rat_18_valid <= 1'b1;
        end
        if(when_RAT_l30_91) begin
          rat_18_valid <= 1'b1;
        end
        if(when_RAT_l30_92) begin
          rat_18_valid <= 1'b1;
        end
        if(when_RAT_l30_93) begin
          rat_18_valid <= 1'b1;
        end
        if(when_RAT_l30_94) begin
          rat_18_valid <= 1'b1;
        end
        if(when_RAT_l30_95) begin
          rat_19_valid <= 1'b1;
        end
        if(when_RAT_l30_96) begin
          rat_19_valid <= 1'b1;
        end
        if(when_RAT_l30_97) begin
          rat_19_valid <= 1'b1;
        end
        if(when_RAT_l30_98) begin
          rat_19_valid <= 1'b1;
        end
        if(when_RAT_l30_99) begin
          rat_19_valid <= 1'b1;
        end
        if(when_RAT_l30_100) begin
          rat_20_valid <= 1'b1;
        end
        if(when_RAT_l30_101) begin
          rat_20_valid <= 1'b1;
        end
        if(when_RAT_l30_102) begin
          rat_20_valid <= 1'b1;
        end
        if(when_RAT_l30_103) begin
          rat_20_valid <= 1'b1;
        end
        if(when_RAT_l30_104) begin
          rat_20_valid <= 1'b1;
        end
        if(when_RAT_l30_105) begin
          rat_21_valid <= 1'b1;
        end
        if(when_RAT_l30_106) begin
          rat_21_valid <= 1'b1;
        end
        if(when_RAT_l30_107) begin
          rat_21_valid <= 1'b1;
        end
        if(when_RAT_l30_108) begin
          rat_21_valid <= 1'b1;
        end
        if(when_RAT_l30_109) begin
          rat_21_valid <= 1'b1;
        end
        if(when_RAT_l30_110) begin
          rat_22_valid <= 1'b1;
        end
        if(when_RAT_l30_111) begin
          rat_22_valid <= 1'b1;
        end
        if(when_RAT_l30_112) begin
          rat_22_valid <= 1'b1;
        end
        if(when_RAT_l30_113) begin
          rat_22_valid <= 1'b1;
        end
        if(when_RAT_l30_114) begin
          rat_22_valid <= 1'b1;
        end
        if(when_RAT_l30_115) begin
          rat_23_valid <= 1'b1;
        end
        if(when_RAT_l30_116) begin
          rat_23_valid <= 1'b1;
        end
        if(when_RAT_l30_117) begin
          rat_23_valid <= 1'b1;
        end
        if(when_RAT_l30_118) begin
          rat_23_valid <= 1'b1;
        end
        if(when_RAT_l30_119) begin
          rat_23_valid <= 1'b1;
        end
        if(when_RAT_l30_120) begin
          rat_24_valid <= 1'b1;
        end
        if(when_RAT_l30_121) begin
          rat_24_valid <= 1'b1;
        end
        if(when_RAT_l30_122) begin
          rat_24_valid <= 1'b1;
        end
        if(when_RAT_l30_123) begin
          rat_24_valid <= 1'b1;
        end
        if(when_RAT_l30_124) begin
          rat_24_valid <= 1'b1;
        end
        if(when_RAT_l30_125) begin
          rat_25_valid <= 1'b1;
        end
        if(when_RAT_l30_126) begin
          rat_25_valid <= 1'b1;
        end
        if(when_RAT_l30_127) begin
          rat_25_valid <= 1'b1;
        end
        if(when_RAT_l30_128) begin
          rat_25_valid <= 1'b1;
        end
        if(when_RAT_l30_129) begin
          rat_25_valid <= 1'b1;
        end
        if(when_RAT_l30_130) begin
          rat_26_valid <= 1'b1;
        end
        if(when_RAT_l30_131) begin
          rat_26_valid <= 1'b1;
        end
        if(when_RAT_l30_132) begin
          rat_26_valid <= 1'b1;
        end
        if(when_RAT_l30_133) begin
          rat_26_valid <= 1'b1;
        end
        if(when_RAT_l30_134) begin
          rat_26_valid <= 1'b1;
        end
        if(when_RAT_l30_135) begin
          rat_27_valid <= 1'b1;
        end
        if(when_RAT_l30_136) begin
          rat_27_valid <= 1'b1;
        end
        if(when_RAT_l30_137) begin
          rat_27_valid <= 1'b1;
        end
        if(when_RAT_l30_138) begin
          rat_27_valid <= 1'b1;
        end
        if(when_RAT_l30_139) begin
          rat_27_valid <= 1'b1;
        end
        if(when_RAT_l30_140) begin
          rat_28_valid <= 1'b1;
        end
        if(when_RAT_l30_141) begin
          rat_28_valid <= 1'b1;
        end
        if(when_RAT_l30_142) begin
          rat_28_valid <= 1'b1;
        end
        if(when_RAT_l30_143) begin
          rat_28_valid <= 1'b1;
        end
        if(when_RAT_l30_144) begin
          rat_28_valid <= 1'b1;
        end
        if(when_RAT_l30_145) begin
          rat_29_valid <= 1'b1;
        end
        if(when_RAT_l30_146) begin
          rat_29_valid <= 1'b1;
        end
        if(when_RAT_l30_147) begin
          rat_29_valid <= 1'b1;
        end
        if(when_RAT_l30_148) begin
          rat_29_valid <= 1'b1;
        end
        if(when_RAT_l30_149) begin
          rat_29_valid <= 1'b1;
        end
        if(when_RAT_l30_150) begin
          rat_30_valid <= 1'b1;
        end
        if(when_RAT_l30_151) begin
          rat_30_valid <= 1'b1;
        end
        if(when_RAT_l30_152) begin
          rat_30_valid <= 1'b1;
        end
        if(when_RAT_l30_153) begin
          rat_30_valid <= 1'b1;
        end
        if(when_RAT_l30_154) begin
          rat_30_valid <= 1'b1;
        end
        if(when_RAT_l30_155) begin
          rat_31_valid <= 1'b1;
        end
        if(when_RAT_l30_156) begin
          rat_31_valid <= 1'b1;
        end
        if(when_RAT_l30_157) begin
          rat_31_valid <= 1'b1;
        end
        if(when_RAT_l30_158) begin
          rat_31_valid <= 1'b1;
        end
        if(when_RAT_l30_159) begin
          rat_31_valid <= 1'b1;
        end
        if(io_writePort_0_wen) begin
          if(_zz_1[0]) begin
            rat_0_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[1]) begin
            rat_1_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[2]) begin
            rat_2_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[3]) begin
            rat_3_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[4]) begin
            rat_4_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[5]) begin
            rat_5_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[6]) begin
            rat_6_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[7]) begin
            rat_7_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[8]) begin
            rat_8_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[9]) begin
            rat_9_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[10]) begin
            rat_10_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[11]) begin
            rat_11_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[12]) begin
            rat_12_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[13]) begin
            rat_13_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[14]) begin
            rat_14_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[15]) begin
            rat_15_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[16]) begin
            rat_16_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[17]) begin
            rat_17_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[18]) begin
            rat_18_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[19]) begin
            rat_19_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[20]) begin
            rat_20_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[21]) begin
            rat_21_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[22]) begin
            rat_22_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[23]) begin
            rat_23_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[24]) begin
            rat_24_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[25]) begin
            rat_25_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[26]) begin
            rat_26_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[27]) begin
            rat_27_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[28]) begin
            rat_28_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[29]) begin
            rat_29_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[30]) begin
            rat_30_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_1[31]) begin
            rat_31_prfIdx <= io_writePort_0_prd;
          end
          if(_zz_2[0]) begin
            rat_0_valid <= 1'b0;
          end
          if(_zz_2[1]) begin
            rat_1_valid <= 1'b0;
          end
          if(_zz_2[2]) begin
            rat_2_valid <= 1'b0;
          end
          if(_zz_2[3]) begin
            rat_3_valid <= 1'b0;
          end
          if(_zz_2[4]) begin
            rat_4_valid <= 1'b0;
          end
          if(_zz_2[5]) begin
            rat_5_valid <= 1'b0;
          end
          if(_zz_2[6]) begin
            rat_6_valid <= 1'b0;
          end
          if(_zz_2[7]) begin
            rat_7_valid <= 1'b0;
          end
          if(_zz_2[8]) begin
            rat_8_valid <= 1'b0;
          end
          if(_zz_2[9]) begin
            rat_9_valid <= 1'b0;
          end
          if(_zz_2[10]) begin
            rat_10_valid <= 1'b0;
          end
          if(_zz_2[11]) begin
            rat_11_valid <= 1'b0;
          end
          if(_zz_2[12]) begin
            rat_12_valid <= 1'b0;
          end
          if(_zz_2[13]) begin
            rat_13_valid <= 1'b0;
          end
          if(_zz_2[14]) begin
            rat_14_valid <= 1'b0;
          end
          if(_zz_2[15]) begin
            rat_15_valid <= 1'b0;
          end
          if(_zz_2[16]) begin
            rat_16_valid <= 1'b0;
          end
          if(_zz_2[17]) begin
            rat_17_valid <= 1'b0;
          end
          if(_zz_2[18]) begin
            rat_18_valid <= 1'b0;
          end
          if(_zz_2[19]) begin
            rat_19_valid <= 1'b0;
          end
          if(_zz_2[20]) begin
            rat_20_valid <= 1'b0;
          end
          if(_zz_2[21]) begin
            rat_21_valid <= 1'b0;
          end
          if(_zz_2[22]) begin
            rat_22_valid <= 1'b0;
          end
          if(_zz_2[23]) begin
            rat_23_valid <= 1'b0;
          end
          if(_zz_2[24]) begin
            rat_24_valid <= 1'b0;
          end
          if(_zz_2[25]) begin
            rat_25_valid <= 1'b0;
          end
          if(_zz_2[26]) begin
            rat_26_valid <= 1'b0;
          end
          if(_zz_2[27]) begin
            rat_27_valid <= 1'b0;
          end
          if(_zz_2[28]) begin
            rat_28_valid <= 1'b0;
          end
          if(_zz_2[29]) begin
            rat_29_valid <= 1'b0;
          end
          if(_zz_2[30]) begin
            rat_30_valid <= 1'b0;
          end
          if(_zz_2[31]) begin
            rat_31_valid <= 1'b0;
          end
        end
        if(io_writePort_1_wen) begin
          if(_zz_3[0]) begin
            rat_0_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[1]) begin
            rat_1_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[2]) begin
            rat_2_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[3]) begin
            rat_3_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[4]) begin
            rat_4_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[5]) begin
            rat_5_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[6]) begin
            rat_6_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[7]) begin
            rat_7_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[8]) begin
            rat_8_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[9]) begin
            rat_9_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[10]) begin
            rat_10_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[11]) begin
            rat_11_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[12]) begin
            rat_12_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[13]) begin
            rat_13_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[14]) begin
            rat_14_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[15]) begin
            rat_15_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[16]) begin
            rat_16_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[17]) begin
            rat_17_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[18]) begin
            rat_18_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[19]) begin
            rat_19_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[20]) begin
            rat_20_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[21]) begin
            rat_21_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[22]) begin
            rat_22_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[23]) begin
            rat_23_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[24]) begin
            rat_24_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[25]) begin
            rat_25_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[26]) begin
            rat_26_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[27]) begin
            rat_27_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[28]) begin
            rat_28_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[29]) begin
            rat_29_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[30]) begin
            rat_30_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_3[31]) begin
            rat_31_prfIdx <= io_writePort_1_prd;
          end
          if(_zz_4[0]) begin
            rat_0_valid <= 1'b0;
          end
          if(_zz_4[1]) begin
            rat_1_valid <= 1'b0;
          end
          if(_zz_4[2]) begin
            rat_2_valid <= 1'b0;
          end
          if(_zz_4[3]) begin
            rat_3_valid <= 1'b0;
          end
          if(_zz_4[4]) begin
            rat_4_valid <= 1'b0;
          end
          if(_zz_4[5]) begin
            rat_5_valid <= 1'b0;
          end
          if(_zz_4[6]) begin
            rat_6_valid <= 1'b0;
          end
          if(_zz_4[7]) begin
            rat_7_valid <= 1'b0;
          end
          if(_zz_4[8]) begin
            rat_8_valid <= 1'b0;
          end
          if(_zz_4[9]) begin
            rat_9_valid <= 1'b0;
          end
          if(_zz_4[10]) begin
            rat_10_valid <= 1'b0;
          end
          if(_zz_4[11]) begin
            rat_11_valid <= 1'b0;
          end
          if(_zz_4[12]) begin
            rat_12_valid <= 1'b0;
          end
          if(_zz_4[13]) begin
            rat_13_valid <= 1'b0;
          end
          if(_zz_4[14]) begin
            rat_14_valid <= 1'b0;
          end
          if(_zz_4[15]) begin
            rat_15_valid <= 1'b0;
          end
          if(_zz_4[16]) begin
            rat_16_valid <= 1'b0;
          end
          if(_zz_4[17]) begin
            rat_17_valid <= 1'b0;
          end
          if(_zz_4[18]) begin
            rat_18_valid <= 1'b0;
          end
          if(_zz_4[19]) begin
            rat_19_valid <= 1'b0;
          end
          if(_zz_4[20]) begin
            rat_20_valid <= 1'b0;
          end
          if(_zz_4[21]) begin
            rat_21_valid <= 1'b0;
          end
          if(_zz_4[22]) begin
            rat_22_valid <= 1'b0;
          end
          if(_zz_4[23]) begin
            rat_23_valid <= 1'b0;
          end
          if(_zz_4[24]) begin
            rat_24_valid <= 1'b0;
          end
          if(_zz_4[25]) begin
            rat_25_valid <= 1'b0;
          end
          if(_zz_4[26]) begin
            rat_26_valid <= 1'b0;
          end
          if(_zz_4[27]) begin
            rat_27_valid <= 1'b0;
          end
          if(_zz_4[28]) begin
            rat_28_valid <= 1'b0;
          end
          if(_zz_4[29]) begin
            rat_29_valid <= 1'b0;
          end
          if(_zz_4[30]) begin
            rat_30_valid <= 1'b0;
          end
          if(_zz_4[31]) begin
            rat_31_valid <= 1'b0;
          end
        end
      end
    end
  end


endmodule

module MemService (
  input  wire          io_input_valid,
  input  wire [3:0]    io_input_payload_uop_lsuOp,
  input  wire [4:0]    io_input_payload_uop_lsuCoOp,
  input  wire [31:0]   io_input_payload_vaddr,
  input  wire [9:0]    io_input_payload_asid,
  input  wire          io_iCacheCtrl_busy,
  output reg           io_iCacheCtrl_stall,
  output wire [31:0]   io_iCacheCtrl_cacopVA,
  output wire          io_iCacheCtrl_cacopStoreTag,
  output wire          io_iCacheCtrl_cacopIndexInvalidate,
  output wire          io_iCacheCtrl_cacopHitInvalidate,
  input  wire          io_dCacheCtrl_busy,
  output reg           io_dCacheCtrl_stall,
  output wire [31:0]   io_dCacheCtrl_cacopVA,
  output wire          io_dCacheCtrl_cacopStoreTag,
  output wire          io_dCacheCtrl_cacopIndexInvalidate,
  output wire          io_dCacheCtrl_cacopHitInvalidate,
  output wire [2:0]    io_TLBCtrl_op,
  output wire          io_TLBCtrl_invGlobal,
  output wire          io_TLBCtrl_invLocal,
  output wire          io_TLBCtrl_invLocalVAMatch,
  output wire          io_TLBCtrl_invLocalVANotMatch,
  output wire [1:0]    io_TLBCtrl_index,
  output wire [18:0]   io_TLBCtrl_invVA,
  output wire [9:0]    io_TLBCtrl_asid,
  input  wire          io_flush,
  input  wire          io_wake,
  input  wire          aclk,
  input  wire          aresetn
);
  localparam LSUOp_cacop = 4'd0;
  localparam LSUOp_tlbsrch = 4'd1;
  localparam LSUOp_tlbrd = 4'd2;
  localparam LSUOp_tlbwr = 4'd3;
  localparam LSUOp_tlbfill = 4'd4;
  localparam LSUOp_invtlb = 4'd5;
  localparam LSUOp_ll = 4'd6;
  localparam LSUOp_sc = 4'd7;
  localparam LSUOp_ld = 4'd8;
  localparam LSUOp_ldu = 4'd9;
  localparam LSUOp_st = 4'd10;
  localparam LSUOp_preld = 4'd11;
  localparam LSUOp_dbar = 4'd12;
  localparam LSUOp_ibar = 4'd13;
  localparam TLBOp_nop = 3'd0;
  localparam TLBOp_srch = 3'd1;
  localparam TLBOp_read = 3'd2;
  localparam TLBOp_write = 3'd3;
  localparam TLBOp_fill = 3'd4;
  localparam TLBOp_inv = 3'd5;
  localparam fsm_enumDef_BOOT = 3'd0;
  localparam fsm_enumDef_idle = 3'd1;
  localparam fsm_enumDef_waitToBegin = 3'd2;
  localparam fsm_enumDef_waitToFinish = 3'd3;
  localparam fsm_enumDef_cacop = 3'd4;
  localparam fsm_enumDef_tlb = 3'd5;

  wire       [1:0]    _zz_invCounter_valueNext;
  wire       [0:0]    _zz_invCounter_valueNext_1;
  wire       [1:0]    _zz_iCacheIndexInvalidate;
  wire       [0:0]    _zz_iCacheIndexInvalidate_1;
  wire       [1:0]    _zz_dCacheIndexInvalidate;
  wire       [0:0]    _zz_dCacheIndexInvalidate_1;
  wire       [4:0]    _zz_tlbInvGlobal;
  wire       [0:0]    _zz_tlbInvGlobal_1;
  wire       [4:0]    _zz_tlbInvGlobal_2;
  wire       [1:0]    _zz_tlbInvGlobal_3;
  wire       [4:0]    _zz_tlbInvGlobal_4;
  wire       [2:0]    _zz_tlbInvGlobal_5;
  wire       [4:0]    _zz_tlbInvLocal;
  wire       [0:0]    _zz_tlbInvLocal_1;
  wire       [4:0]    _zz_tlbInvLocal_2;
  wire       [1:0]    _zz_tlbInvLocal_3;
  wire       [4:0]    _zz_tlbInvLocalVAMatch;
  wire       [2:0]    _zz_tlbInvLocalVAMatch_1;
  wire       [4:0]    _zz_tlbInvLocalVAMatch_2;
  wire       [2:0]    _zz_tlbInvLocalVAMatch_3;
  wire       [4:0]    _zz_tlbInvLocalVAMatch_4;
  wire       [2:0]    _zz_tlbInvLocalVAMatch_5;
  wire       [4:0]    _zz_tlbInvLocalVANotMatch;
  wire       [2:0]    _zz_tlbInvLocalVANotMatch_1;
  reg        [3:0]    opBuffer_op;
  reg        [4:0]    opBuffer_hint;
  reg        [31:0]   opBuffer_vaddr;
  reg        [9:0]    opBuffer_asid;
  reg                 bufferLock;
  wire                when_MEMService_l26;
  wire                when_MEMService_l32;
  reg                 iCacheStoreTag;
  reg                 iCacheIndexInvalidate;
  reg                 iCacheHitInvalidate;
  reg                 dCacheStoreTag;
  reg                 dCacheIndexInvalidate;
  reg                 dCacheHitInvalidate;
  reg        [2:0]    tlbOp_1;
  reg                 tlbInvGlobal;
  reg                 tlbInvLocal;
  reg                 tlbInvLocalVAMatch;
  reg                 tlbInvLocalVANotMatch;
  reg                 invCounter_willIncrement;
  reg                 invCounter_willClear;
  reg        [1:0]    invCounter_valueNext;
  reg        [1:0]    invCounter_value;
  wire                invCounter_willOverflowIfInc;
  wire                invCounter_willOverflow;
  reg        [2:0]    tlbOpNext;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg        [2:0]    fsm_stateReg;
  reg        [2:0]    fsm_stateNext;
  wire                when_MEMService_l113;
  wire                when_MEMService_l114;
  wire                when_MEMService_l123;
  wire                when_MEMService_l183;
  wire                when_MEMService_l156;
  wire                when_MEMService_l159;
  `ifndef SYNTHESIS
  reg [55:0] io_input_payload_uop_lsuOp_string;
  reg [39:0] io_TLBCtrl_op_string;
  reg [55:0] opBuffer_op_string;
  reg [39:0] tlbOp_1_string;
  reg [39:0] tlbOpNext_string;
  reg [95:0] fsm_stateReg_string;
  reg [95:0] fsm_stateNext_string;
  `endif


  assign _zz_invCounter_valueNext_1 = invCounter_willIncrement;
  assign _zz_invCounter_valueNext = {1'd0, _zz_invCounter_valueNext_1};
  assign _zz_iCacheIndexInvalidate_1 = 1'b1;
  assign _zz_iCacheIndexInvalidate = {1'd0, _zz_iCacheIndexInvalidate_1};
  assign _zz_dCacheIndexInvalidate_1 = 1'b1;
  assign _zz_dCacheIndexInvalidate = {1'd0, _zz_dCacheIndexInvalidate_1};
  assign _zz_tlbInvGlobal_1 = 1'b1;
  assign _zz_tlbInvGlobal = {4'd0, _zz_tlbInvGlobal_1};
  assign _zz_tlbInvGlobal_3 = 2'b10;
  assign _zz_tlbInvGlobal_2 = {3'd0, _zz_tlbInvGlobal_3};
  assign _zz_tlbInvGlobal_5 = 3'b110;
  assign _zz_tlbInvGlobal_4 = {2'd0, _zz_tlbInvGlobal_5};
  assign _zz_tlbInvLocal_1 = 1'b1;
  assign _zz_tlbInvLocal = {4'd0, _zz_tlbInvLocal_1};
  assign _zz_tlbInvLocal_3 = 2'b11;
  assign _zz_tlbInvLocal_2 = {3'd0, _zz_tlbInvLocal_3};
  assign _zz_tlbInvLocalVAMatch_1 = 3'b100;
  assign _zz_tlbInvLocalVAMatch = {2'd0, _zz_tlbInvLocalVAMatch_1};
  assign _zz_tlbInvLocalVAMatch_3 = 3'b101;
  assign _zz_tlbInvLocalVAMatch_2 = {2'd0, _zz_tlbInvLocalVAMatch_3};
  assign _zz_tlbInvLocalVAMatch_5 = 3'b110;
  assign _zz_tlbInvLocalVAMatch_4 = {2'd0, _zz_tlbInvLocalVAMatch_5};
  assign _zz_tlbInvLocalVANotMatch_1 = 3'b100;
  assign _zz_tlbInvLocalVANotMatch = {2'd0, _zz_tlbInvLocalVANotMatch_1};
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_uop_lsuOp)
      LSUOp_cacop : io_input_payload_uop_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : io_input_payload_uop_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : io_input_payload_uop_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : io_input_payload_uop_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : io_input_payload_uop_lsuOp_string = "tlbfill";
      LSUOp_invtlb : io_input_payload_uop_lsuOp_string = "invtlb ";
      LSUOp_ll : io_input_payload_uop_lsuOp_string = "ll     ";
      LSUOp_sc : io_input_payload_uop_lsuOp_string = "sc     ";
      LSUOp_ld : io_input_payload_uop_lsuOp_string = "ld     ";
      LSUOp_ldu : io_input_payload_uop_lsuOp_string = "ldu    ";
      LSUOp_st : io_input_payload_uop_lsuOp_string = "st     ";
      LSUOp_preld : io_input_payload_uop_lsuOp_string = "preld  ";
      LSUOp_dbar : io_input_payload_uop_lsuOp_string = "dbar   ";
      LSUOp_ibar : io_input_payload_uop_lsuOp_string = "ibar   ";
      default : io_input_payload_uop_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_TLBCtrl_op)
      TLBOp_nop : io_TLBCtrl_op_string = "nop  ";
      TLBOp_srch : io_TLBCtrl_op_string = "srch ";
      TLBOp_read : io_TLBCtrl_op_string = "read ";
      TLBOp_write : io_TLBCtrl_op_string = "write";
      TLBOp_fill : io_TLBCtrl_op_string = "fill ";
      TLBOp_inv : io_TLBCtrl_op_string = "inv  ";
      default : io_TLBCtrl_op_string = "?????";
    endcase
  end
  always @(*) begin
    case(opBuffer_op)
      LSUOp_cacop : opBuffer_op_string = "cacop  ";
      LSUOp_tlbsrch : opBuffer_op_string = "tlbsrch";
      LSUOp_tlbrd : opBuffer_op_string = "tlbrd  ";
      LSUOp_tlbwr : opBuffer_op_string = "tlbwr  ";
      LSUOp_tlbfill : opBuffer_op_string = "tlbfill";
      LSUOp_invtlb : opBuffer_op_string = "invtlb ";
      LSUOp_ll : opBuffer_op_string = "ll     ";
      LSUOp_sc : opBuffer_op_string = "sc     ";
      LSUOp_ld : opBuffer_op_string = "ld     ";
      LSUOp_ldu : opBuffer_op_string = "ldu    ";
      LSUOp_st : opBuffer_op_string = "st     ";
      LSUOp_preld : opBuffer_op_string = "preld  ";
      LSUOp_dbar : opBuffer_op_string = "dbar   ";
      LSUOp_ibar : opBuffer_op_string = "ibar   ";
      default : opBuffer_op_string = "???????";
    endcase
  end
  always @(*) begin
    case(tlbOp_1)
      TLBOp_nop : tlbOp_1_string = "nop  ";
      TLBOp_srch : tlbOp_1_string = "srch ";
      TLBOp_read : tlbOp_1_string = "read ";
      TLBOp_write : tlbOp_1_string = "write";
      TLBOp_fill : tlbOp_1_string = "fill ";
      TLBOp_inv : tlbOp_1_string = "inv  ";
      default : tlbOp_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(tlbOpNext)
      TLBOp_nop : tlbOpNext_string = "nop  ";
      TLBOp_srch : tlbOpNext_string = "srch ";
      TLBOp_read : tlbOpNext_string = "read ";
      TLBOp_write : tlbOpNext_string = "write";
      TLBOp_fill : tlbOpNext_string = "fill ";
      TLBOp_inv : tlbOpNext_string = "inv  ";
      default : tlbOpNext_string = "?????";
    endcase
  end
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_BOOT : fsm_stateReg_string = "BOOT        ";
      fsm_enumDef_idle : fsm_stateReg_string = "idle        ";
      fsm_enumDef_waitToBegin : fsm_stateReg_string = "waitToBegin ";
      fsm_enumDef_waitToFinish : fsm_stateReg_string = "waitToFinish";
      fsm_enumDef_cacop : fsm_stateReg_string = "cacop       ";
      fsm_enumDef_tlb : fsm_stateReg_string = "tlb         ";
      default : fsm_stateReg_string = "????????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_BOOT : fsm_stateNext_string = "BOOT        ";
      fsm_enumDef_idle : fsm_stateNext_string = "idle        ";
      fsm_enumDef_waitToBegin : fsm_stateNext_string = "waitToBegin ";
      fsm_enumDef_waitToFinish : fsm_stateNext_string = "waitToFinish";
      fsm_enumDef_cacop : fsm_stateNext_string = "cacop       ";
      fsm_enumDef_tlb : fsm_stateNext_string = "tlb         ";
      default : fsm_stateNext_string = "????????????";
    endcase
  end
  `endif

  assign when_MEMService_l26 = (io_input_valid && (! bufferLock));
  assign when_MEMService_l32 = (io_input_valid && (! io_flush));
  always @(*) begin
    io_iCacheCtrl_stall = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_idle : begin
      end
      fsm_enumDef_waitToBegin : begin
        io_iCacheCtrl_stall = 1'b1;
      end
      fsm_enumDef_waitToFinish : begin
        io_iCacheCtrl_stall = 1'b1;
      end
      fsm_enumDef_cacop : begin
        io_iCacheCtrl_stall = 1'b1;
      end
      fsm_enumDef_tlb : begin
        io_iCacheCtrl_stall = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign io_iCacheCtrl_cacopVA = opBuffer_vaddr;
  assign io_iCacheCtrl_cacopStoreTag = iCacheStoreTag;
  assign io_iCacheCtrl_cacopIndexInvalidate = iCacheIndexInvalidate;
  assign io_iCacheCtrl_cacopHitInvalidate = iCacheHitInvalidate;
  always @(*) begin
    io_dCacheCtrl_stall = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_idle : begin
      end
      fsm_enumDef_waitToBegin : begin
        io_dCacheCtrl_stall = 1'b1;
      end
      fsm_enumDef_waitToFinish : begin
        io_dCacheCtrl_stall = 1'b1;
      end
      fsm_enumDef_cacop : begin
        io_dCacheCtrl_stall = 1'b1;
      end
      fsm_enumDef_tlb : begin
        io_dCacheCtrl_stall = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign io_dCacheCtrl_cacopVA = opBuffer_vaddr;
  assign io_dCacheCtrl_cacopStoreTag = dCacheStoreTag;
  assign io_dCacheCtrl_cacopIndexInvalidate = dCacheIndexInvalidate;
  assign io_dCacheCtrl_cacopHitInvalidate = dCacheHitInvalidate;
  assign io_TLBCtrl_op = tlbOp_1;
  assign io_TLBCtrl_invGlobal = tlbInvGlobal;
  assign io_TLBCtrl_invLocal = tlbInvLocal;
  assign io_TLBCtrl_invLocalVAMatch = tlbInvLocalVAMatch;
  assign io_TLBCtrl_invLocalVANotMatch = tlbInvLocalVANotMatch;
  assign io_TLBCtrl_invVA = opBuffer_vaddr[31 : 13];
  assign io_TLBCtrl_asid = opBuffer_asid;
  always @(*) begin
    invCounter_willIncrement = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_idle : begin
      end
      fsm_enumDef_waitToBegin : begin
      end
      fsm_enumDef_waitToFinish : begin
      end
      fsm_enumDef_cacop : begin
      end
      fsm_enumDef_tlb : begin
        if(when_MEMService_l156) begin
          invCounter_willIncrement = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    invCounter_willClear = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_idle : begin
      end
      fsm_enumDef_waitToBegin : begin
        if(when_MEMService_l113) begin
          if(!when_MEMService_l114) begin
            if(when_MEMService_l123) begin
              invCounter_willClear = 1'b1;
            end
          end
        end
      end
      fsm_enumDef_waitToFinish : begin
      end
      fsm_enumDef_cacop : begin
      end
      fsm_enumDef_tlb : begin
      end
      default : begin
      end
    endcase
  end

  assign invCounter_willOverflowIfInc = (invCounter_value == 2'b11);
  assign invCounter_willOverflow = (invCounter_willOverflowIfInc && invCounter_willIncrement);
  always @(*) begin
    invCounter_valueNext = (invCounter_value + _zz_invCounter_valueNext);
    if(invCounter_willClear) begin
      invCounter_valueNext = 2'b00;
    end
  end

  assign io_TLBCtrl_index = invCounter_value;
  always @(*) begin
    case(opBuffer_op)
      LSUOp_tlbsrch : begin
        tlbOpNext = TLBOp_srch;
      end
      LSUOp_tlbrd : begin
        tlbOpNext = TLBOp_read;
      end
      LSUOp_tlbwr : begin
        tlbOpNext = TLBOp_write;
      end
      LSUOp_tlbfill : begin
        tlbOpNext = TLBOp_fill;
      end
      LSUOp_invtlb : begin
        tlbOpNext = TLBOp_inv;
      end
      default : begin
        tlbOpNext = TLBOp_nop;
      end
    endcase
  end

  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_idle : begin
      end
      fsm_enumDef_waitToBegin : begin
      end
      fsm_enumDef_waitToFinish : begin
      end
      fsm_enumDef_cacop : begin
      end
      fsm_enumDef_tlb : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_enumDef_idle : begin
        if(io_wake) begin
          fsm_stateNext = fsm_enumDef_waitToBegin;
        end
      end
      fsm_enumDef_waitToBegin : begin
        if(when_MEMService_l113) begin
          if(when_MEMService_l114) begin
            fsm_stateNext = fsm_enumDef_cacop;
          end else begin
            if(when_MEMService_l123) begin
              fsm_stateNext = fsm_enumDef_tlb;
            end else begin
              fsm_stateNext = fsm_enumDef_idle;
            end
          end
        end
      end
      fsm_enumDef_waitToFinish : begin
        if(when_MEMService_l183) begin
          fsm_stateNext = fsm_enumDef_idle;
        end
      end
      fsm_enumDef_cacop : begin
        fsm_stateNext = fsm_enumDef_waitToFinish;
      end
      fsm_enumDef_tlb : begin
        if(when_MEMService_l156) begin
          if(when_MEMService_l159) begin
            fsm_stateNext = fsm_enumDef_idle;
          end
        end else begin
          fsm_stateNext = fsm_enumDef_idle;
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_enumDef_idle;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_BOOT;
    end
  end

  assign when_MEMService_l113 = (! (io_iCacheCtrl_busy || io_dCacheCtrl_busy));
  assign when_MEMService_l114 = (opBuffer_op == LSUOp_cacop);
  assign when_MEMService_l123 = ((((opBuffer_op == LSUOp_tlbsrch) || (opBuffer_op == LSUOp_tlbwr)) || (opBuffer_op == LSUOp_tlbfill)) || (opBuffer_op == LSUOp_invtlb));
  assign when_MEMService_l183 = (! (io_iCacheCtrl_busy || io_dCacheCtrl_busy));
  assign when_MEMService_l156 = (tlbOp_1 == TLBOp_inv);
  assign when_MEMService_l159 = (invCounter_valueNext == 2'b11);
  always @(posedge aclk) begin
    if(!aresetn) begin
      opBuffer_op <= LSUOp_preld;
      opBuffer_hint <= 5'h00;
      opBuffer_vaddr <= 32'h00000000;
      opBuffer_asid <= 10'h000;
      bufferLock <= 1'b0;
      iCacheStoreTag <= 1'b0;
      iCacheIndexInvalidate <= 1'b0;
      iCacheHitInvalidate <= 1'b0;
      dCacheStoreTag <= 1'b0;
      dCacheIndexInvalidate <= 1'b0;
      dCacheHitInvalidate <= 1'b0;
      tlbOp_1 <= TLBOp_nop;
      tlbInvGlobal <= 1'b0;
      tlbInvLocal <= 1'b0;
      tlbInvLocalVAMatch <= 1'b0;
      tlbInvLocalVANotMatch <= 1'b0;
      invCounter_value <= 2'b00;
      fsm_stateReg <= fsm_enumDef_BOOT;
    end else begin
      if(when_MEMService_l26) begin
        opBuffer_op <= io_input_payload_uop_lsuOp;
        opBuffer_hint <= io_input_payload_uop_lsuCoOp;
        opBuffer_vaddr <= io_input_payload_vaddr;
        opBuffer_asid <= io_input_payload_asid;
      end
      if(when_MEMService_l32) begin
        bufferLock <= 1'b1;
      end
      if(io_flush) begin
        bufferLock <= 1'b0;
      end
      invCounter_value <= invCounter_valueNext;
      fsm_stateReg <= fsm_stateNext;
      case(fsm_stateReg)
        fsm_enumDef_idle : begin
        end
        fsm_enumDef_waitToBegin : begin
          if(when_MEMService_l113) begin
            if(when_MEMService_l114) begin
              iCacheStoreTag <= ((opBuffer_hint[4 : 3] == 2'b00) && (opBuffer_hint[2 : 0] == 3'b000));
              iCacheIndexInvalidate <= ((opBuffer_hint[4 : 3] == _zz_iCacheIndexInvalidate) && (opBuffer_hint[2 : 0] == 3'b000));
              iCacheHitInvalidate <= ((opBuffer_hint[4 : 3] == 2'b10) && (opBuffer_hint[2 : 0] == 3'b000));
              dCacheStoreTag <= ((opBuffer_hint[4 : 3] == 2'b00) && (! (opBuffer_hint[2 : 0] == 3'b000)));
              dCacheIndexInvalidate <= ((opBuffer_hint[4 : 3] == _zz_dCacheIndexInvalidate) && (! (opBuffer_hint[2 : 0] == 3'b000)));
              dCacheHitInvalidate <= ((opBuffer_hint[4 : 3] == 2'b10) && (! (opBuffer_hint[2 : 0] == 3'b000)));
            end else begin
              if(when_MEMService_l123) begin
                tlbOp_1 <= tlbOpNext;
                tlbInvGlobal <= ((((opBuffer_hint == 5'h00) || (opBuffer_hint == _zz_tlbInvGlobal)) || (opBuffer_hint == _zz_tlbInvGlobal_2)) || (opBuffer_hint == _zz_tlbInvGlobal_4));
                tlbInvLocal <= (((opBuffer_hint == 5'h00) || (opBuffer_hint == _zz_tlbInvLocal)) || (opBuffer_hint == _zz_tlbInvLocal_2));
                tlbInvLocalVAMatch <= (((opBuffer_hint == _zz_tlbInvLocalVAMatch) || (opBuffer_hint == _zz_tlbInvLocalVAMatch_2)) || (opBuffer_hint == _zz_tlbInvLocalVAMatch_4));
                tlbInvLocalVANotMatch <= (opBuffer_hint == _zz_tlbInvLocalVANotMatch);
              end
            end
          end
        end
        fsm_enumDef_waitToFinish : begin
        end
        fsm_enumDef_cacop : begin
          iCacheStoreTag <= 1'b0;
          iCacheIndexInvalidate <= 1'b0;
          iCacheHitInvalidate <= 1'b0;
          dCacheStoreTag <= 1'b0;
          dCacheIndexInvalidate <= 1'b0;
          dCacheHitInvalidate <= 1'b0;
        end
        fsm_enumDef_tlb : begin
          if(when_MEMService_l156) begin
            if(when_MEMService_l159) begin
              tlbOp_1 <= TLBOp_nop;
              tlbInvGlobal <= 1'b0;
              tlbInvLocal <= 1'b0;
              tlbInvLocalVAMatch <= 1'b0;
              tlbInvLocalVANotMatch <= 1'b0;
            end
          end else begin
            tlbOp_1 <= TLBOp_nop;
            tlbInvGlobal <= 1'b0;
            tlbInvLocal <= 1'b0;
            tlbInvLocalVAMatch <= 1'b0;
            tlbInvLocalVANotMatch <= 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end


endmodule

module TLB (
  output reg           io_iCacheReq_hit,
  output reg  [19:0]   io_iCacheReq_pageInfo_ppn,
  output reg  [1:0]    io_iCacheReq_pageInfo_plv,
  output reg  [1:0]    io_iCacheReq_pageInfo_mat,
  output reg           io_iCacheReq_pageInfo_d,
  output reg           io_iCacheReq_pageInfo_v,
  input  wire [19:0]   io_iCacheReq_virtPageNumber,
  output reg           io_dCacheReq_hit,
  output reg  [19:0]   io_dCacheReq_pageInfo_ppn,
  output reg  [1:0]    io_dCacheReq_pageInfo_plv,
  output reg  [1:0]    io_dCacheReq_pageInfo_mat,
  output reg           io_dCacheReq_pageInfo_d,
  output reg           io_dCacheReq_pageInfo_v,
  input  wire [19:0]   io_dCacheReq_virtPageNumber,
  input  wire [9:0]    io_csrInfo_asid,
  input  wire [1:0]    _zz_io_iCacheReq_pageInfo_plv,
  input  wire          _zz_when_TLB_l177,
  input  wire          _zz_when_TLB_l177_1,
  input  wire [1:0]    _zz_io_iCacheReq_pageInfo_mat,
  input  wire [1:0]    _zz_io_dCacheReq_pageInfo_mat,
  input  wire          _zz_when_TLB_l178,
  input  wire          _zz_when_TLB_l178_1,
  input  wire [1:0]    _zz_io_iCacheReq_pageInfo_mat_1,
  input  wire [2:0]    _zz_io_iCacheReq_pageInfo_ppn,
  input  wire [2:0]    _zz_when_TLB_l178_2,
  input  wire          _zz_when_TLB_l185,
  input  wire          _zz_when_TLB_l185_1,
  input  wire [1:0]    _zz_io_iCacheReq_pageInfo_mat_2,
  input  wire [2:0]    _zz_io_iCacheReq_pageInfo_ppn_1,
  input  wire [2:0]    _zz_when_TLB_l185_2,
  input  wire [5:0]    _zz_entryToFill_e,
  input  wire [1:0]    _zz_io_csrWrite_asid,
  input  wire [21:0]   _zz_io_swRead_value,
  input  wire [5:0]    _zz_entryToFill_ps,
  input  wire          _zz_io_swRead_value_1,
  input  wire          _zz_entryToFill_e_1,
  input  wire [18:0]   _zz_entryToFill_vppn,
  input  wire          _zz_entryToFill_pp0_v,
  input  wire          _zz_entryToFill_pp0_d,
  input  wire [1:0]    _zz_entryToFill_pp0_plv,
  input  wire [1:0]    _zz_entryToFill_pp0_mat,
  input  wire          _zz_entryToFill_g,
  input  wire [19:0]   _zz_entryToFill_pp0_ppn,
  input  wire          _zz_entryToFill_pp1_v,
  input  wire          _zz_entryToFill_pp1_d,
  input  wire [1:0]    _zz_entryToFill_pp1_plv,
  input  wire [1:0]    _zz_entryToFill_pp1_mat,
  input  wire          _zz_entryToFill_g_1,
  input  wire [19:0]   _zz_entryToFill_pp1_ppn,
  output reg  [1:0]    _zz_io_swRead_value_2,
  output reg  [21:0]   _zz_io_swRead_value_3,
  output reg  [5:0]    _zz_io_swRead_value_4,
  output reg           _zz_io_swRead_value_5,
  output reg           _zz_io_swRead_value_6,
  output reg  [12:0]   _zz_io_swRead_value_7,
  output reg  [18:0]   _zz_io_swRead_value_8,
  output reg           _zz_io_swRead_value_9,
  output reg           _zz_io_swRead_value_10,
  output reg  [1:0]    _zz_io_swRead_value_11,
  output reg  [1:0]    _zz_io_swRead_value_12,
  output reg           _zz_io_swRead_value_13,
  output reg           _zz_io_swRead_value_14,
  output reg  [19:0]   _zz_io_swRead_value_15,
  output reg  [3:0]    _zz_io_swRead_value_16,
  output reg           _zz_io_swRead_value_17,
  output reg           _zz_io_swRead_value_18,
  output reg  [1:0]    _zz_io_swRead_value_19,
  output reg  [1:0]    _zz_io_swRead_value_20,
  output reg           _zz_io_swRead_value_21,
  output reg           _zz_io_swRead_value_22,
  output reg  [19:0]   _zz_io_swRead_value_23,
  output reg  [3:0]    _zz_io_swRead_value_24,
  output reg  [9:0]    io_csrWrite_asid,
  output reg           io_csrWrite_idxWen,
  output reg           io_csrWrite_entryWen,
  input  wire [2:0]    io_ctrl_op,
  input  wire          io_ctrl_invGlobal,
  input  wire          io_ctrl_invLocal,
  input  wire          io_ctrl_invLocalVAMatch,
  input  wire          io_ctrl_invLocalVANotMatch,
  input  wire [1:0]    io_ctrl_index,
  input  wire [18:0]   io_ctrl_invVA,
  input  wire [9:0]    io_ctrl_asid,
  input  wire          aclk,
  input  wire          aresetn
);
  localparam TLBOp_nop = 3'd0;
  localparam TLBOp_srch = 3'd1;
  localparam TLBOp_read = 3'd2;
  localparam TLBOp_write = 3'd3;
  localparam TLBOp_fill = 3'd4;
  localparam TLBOp_inv = 3'd5;

  reg        [19:0]   _zz__zz_io_iCacheReq_pageInfo_ppn_5;
  reg                 _zz__zz_io_iCacheReq_pageInfo_ppn_6;
  reg        [19:0]   _zz_io_iCacheReq_pageInfo_ppn_7;
  reg        [19:0]   _zz_io_iCacheReq_pageInfo_ppn_8;
  reg        [1:0]    _zz_io_iCacheReq_pageInfo_plv_1;
  reg        [1:0]    _zz_io_iCacheReq_pageInfo_plv_2;
  reg        [1:0]    _zz_io_iCacheReq_pageInfo_mat_3;
  reg        [1:0]    _zz_io_iCacheReq_pageInfo_mat_4;
  reg                 _zz_io_iCacheReq_pageInfo_d;
  reg                 _zz_io_iCacheReq_pageInfo_d_1;
  reg                 _zz_io_iCacheReq_pageInfo_v;
  reg                 _zz_io_iCacheReq_pageInfo_v_1;
  reg        [19:0]   _zz__zz_io_dCacheReq_pageInfo_ppn_3;
  reg                 _zz__zz_io_dCacheReq_pageInfo_ppn_4;
  reg        [19:0]   _zz_io_dCacheReq_pageInfo_ppn_5;
  reg        [19:0]   _zz_io_dCacheReq_pageInfo_ppn_6;
  reg        [1:0]    _zz_io_dCacheReq_pageInfo_plv;
  reg        [1:0]    _zz_io_dCacheReq_pageInfo_plv_1;
  reg        [1:0]    _zz_io_dCacheReq_pageInfo_mat_1;
  reg        [1:0]    _zz_io_dCacheReq_pageInfo_mat_2;
  reg                 _zz_io_dCacheReq_pageInfo_d;
  reg                 _zz_io_dCacheReq_pageInfo_d_1;
  reg                 _zz_io_dCacheReq_pageInfo_v;
  reg                 _zz_io_dCacheReq_pageInfo_v_1;
  wire       [1:0]    _zz_replaceCounter_valueNext;
  wire       [0:0]    _zz_replaceCounter_valueNext_1;
  reg                 _zz__zz_io_csrWrite_asid_1;
  wire       [1:0]    _zz__zz_io_csrWrite_asid_1_1;
  reg        [5:0]    _zz__zz_io_swRead_value_4;
  wire       [1:0]    _zz__zz_io_swRead_value_4_1;
  reg        [18:0]   _zz__zz_io_swRead_value_8;
  wire       [1:0]    _zz__zz_io_swRead_value_8_1;
  reg                 _zz__zz_io_swRead_value_9;
  wire       [1:0]    _zz__zz_io_swRead_value_9_1;
  reg                 _zz__zz_io_swRead_value_10;
  wire       [1:0]    _zz__zz_io_swRead_value_10_1;
  reg        [1:0]    _zz__zz_io_swRead_value_11;
  wire       [1:0]    _zz__zz_io_swRead_value_11_1;
  reg        [1:0]    _zz__zz_io_swRead_value_12;
  wire       [1:0]    _zz__zz_io_swRead_value_12_1;
  reg                 _zz__zz_io_swRead_value_13;
  wire       [1:0]    _zz__zz_io_swRead_value_13_1;
  reg        [19:0]   _zz__zz_io_swRead_value_15;
  wire       [1:0]    _zz__zz_io_swRead_value_15_1;
  reg                 _zz__zz_io_swRead_value_17;
  wire       [1:0]    _zz__zz_io_swRead_value_17_1;
  reg                 _zz__zz_io_swRead_value_18;
  wire       [1:0]    _zz__zz_io_swRead_value_18_1;
  reg        [1:0]    _zz__zz_io_swRead_value_19;
  wire       [1:0]    _zz__zz_io_swRead_value_19_1;
  reg        [1:0]    _zz__zz_io_swRead_value_20;
  wire       [1:0]    _zz__zz_io_swRead_value_20_1;
  reg                 _zz__zz_io_swRead_value_21;
  wire       [1:0]    _zz__zz_io_swRead_value_21_1;
  reg        [19:0]   _zz__zz_io_swRead_value_23;
  wire       [1:0]    _zz__zz_io_swRead_value_23_1;
  reg                 _zz__zz_when_TLB_l130;
  reg        [9:0]    _zz__zz_when_TLB_l130_1;
  reg        [18:0]   _zz__zz_when_TLB_l130_2;
  wire       [19:0]   _zz__zz_when_TLB_l130_2_1;
  reg        [5:0]    _zz__zz_when_TLB_l130_2_2;
  reg        [18:0]   tlbStorage_0_vppn;
  reg        [5:0]    tlbStorage_0_ps;
  reg                 tlbStorage_0_g;
  reg        [9:0]    tlbStorage_0_asid;
  reg                 tlbStorage_0_e;
  reg        [19:0]   tlbStorage_0_pp0_ppn;
  reg        [1:0]    tlbStorage_0_pp0_plv;
  reg        [1:0]    tlbStorage_0_pp0_mat;
  reg                 tlbStorage_0_pp0_d;
  reg                 tlbStorage_0_pp0_v;
  reg        [19:0]   tlbStorage_0_pp1_ppn;
  reg        [1:0]    tlbStorage_0_pp1_plv;
  reg        [1:0]    tlbStorage_0_pp1_mat;
  reg                 tlbStorage_0_pp1_d;
  reg                 tlbStorage_0_pp1_v;
  reg        [18:0]   tlbStorage_1_vppn;
  reg        [5:0]    tlbStorage_1_ps;
  reg                 tlbStorage_1_g;
  reg        [9:0]    tlbStorage_1_asid;
  reg                 tlbStorage_1_e;
  reg        [19:0]   tlbStorage_1_pp0_ppn;
  reg        [1:0]    tlbStorage_1_pp0_plv;
  reg        [1:0]    tlbStorage_1_pp0_mat;
  reg                 tlbStorage_1_pp0_d;
  reg                 tlbStorage_1_pp0_v;
  reg        [19:0]   tlbStorage_1_pp1_ppn;
  reg        [1:0]    tlbStorage_1_pp1_plv;
  reg        [1:0]    tlbStorage_1_pp1_mat;
  reg                 tlbStorage_1_pp1_d;
  reg                 tlbStorage_1_pp1_v;
  reg        [18:0]   tlbStorage_2_vppn;
  reg        [5:0]    tlbStorage_2_ps;
  reg                 tlbStorage_2_g;
  reg        [9:0]    tlbStorage_2_asid;
  reg                 tlbStorage_2_e;
  reg        [19:0]   tlbStorage_2_pp0_ppn;
  reg        [1:0]    tlbStorage_2_pp0_plv;
  reg        [1:0]    tlbStorage_2_pp0_mat;
  reg                 tlbStorage_2_pp0_d;
  reg                 tlbStorage_2_pp0_v;
  reg        [19:0]   tlbStorage_2_pp1_ppn;
  reg        [1:0]    tlbStorage_2_pp1_plv;
  reg        [1:0]    tlbStorage_2_pp1_mat;
  reg                 tlbStorage_2_pp1_d;
  reg                 tlbStorage_2_pp1_v;
  reg        [18:0]   tlbStorage_3_vppn;
  reg        [5:0]    tlbStorage_3_ps;
  reg                 tlbStorage_3_g;
  reg        [9:0]    tlbStorage_3_asid;
  reg                 tlbStorage_3_e;
  reg        [19:0]   tlbStorage_3_pp0_ppn;
  reg        [1:0]    tlbStorage_3_pp0_plv;
  reg        [1:0]    tlbStorage_3_pp0_mat;
  reg                 tlbStorage_3_pp0_d;
  reg                 tlbStorage_3_pp0_v;
  reg        [19:0]   tlbStorage_3_pp1_ppn;
  reg        [1:0]    tlbStorage_3_pp1_plv;
  reg        [1:0]    tlbStorage_3_pp1_mat;
  reg                 tlbStorage_3_pp1_d;
  reg                 tlbStorage_3_pp1_v;
  wire                when_TLB_l177;
  wire                when_TLB_l178;
  wire                _zz_io_iCacheReq_hit;
  wire                _zz_io_iCacheReq_hit_1;
  wire                _zz_io_iCacheReq_hit_2;
  wire       [19:0]   _zz_io_iCacheReq_hit_3;
  wire       [19:0]   _zz_io_iCacheReq_hit_4;
  wire       [19:0]   _zz_io_iCacheReq_hit_5;
  wire       [19:0]   _zz_io_iCacheReq_hit_6;
  wire                _zz_io_iCacheReq_pageInfo_ppn_2;
  wire                _zz_io_iCacheReq_pageInfo_ppn_3;
  wire       [1:0]    _zz_io_iCacheReq_pageInfo_ppn_4;
  wire       [19:0]   _zz_io_iCacheReq_pageInfo_ppn_5;
  wire                _zz_io_iCacheReq_pageInfo_ppn_6;
  wire                _zz_io_iCacheReq_hit_7;
  wire                when_TLB_l185;
  wire                when_TLB_l195;
  wire                when_TLB_l177_1;
  wire                when_TLB_l178_1;
  wire                _zz_io_dCacheReq_hit;
  wire                _zz_io_dCacheReq_hit_1;
  wire                _zz_io_dCacheReq_hit_2;
  wire       [19:0]   _zz_io_dCacheReq_hit_3;
  wire       [19:0]   _zz_io_dCacheReq_hit_4;
  wire       [19:0]   _zz_io_dCacheReq_hit_5;
  wire       [19:0]   _zz_io_dCacheReq_hit_6;
  wire                _zz_io_dCacheReq_pageInfo_ppn;
  wire                _zz_io_dCacheReq_pageInfo_ppn_1;
  wire       [1:0]    _zz_io_dCacheReq_pageInfo_ppn_2;
  wire       [19:0]   _zz_io_dCacheReq_pageInfo_ppn_3;
  wire                _zz_io_dCacheReq_pageInfo_ppn_4;
  wire                _zz_io_dCacheReq_hit_7;
  wire                when_TLB_l185_1;
  wire                when_TLB_l195_1;
  wire       [18:0]   entryToFill_vppn;
  wire       [5:0]    entryToFill_ps;
  wire                entryToFill_g;
  wire       [9:0]    entryToFill_asid;
  wire                entryToFill_e;
  wire       [19:0]   entryToFill_pp0_ppn;
  wire       [1:0]    entryToFill_pp0_plv;
  wire       [1:0]    entryToFill_pp0_mat;
  wire                entryToFill_pp0_d;
  wire                entryToFill_pp0_v;
  wire       [19:0]   entryToFill_pp1_ppn;
  wire       [1:0]    entryToFill_pp1_plv;
  wire       [1:0]    entryToFill_pp1_mat;
  wire                entryToFill_pp1_d;
  wire                entryToFill_pp1_v;
  reg                 replaceCounter_willIncrement;
  wire                replaceCounter_willClear;
  reg        [1:0]    replaceCounter_valueNext;
  reg        [1:0]    replaceCounter_value;
  wire                replaceCounter_willOverflowIfInc;
  wire                replaceCounter_willOverflow;
  wire                _zz_io_swRead_value_25;
  wire                _zz_io_swRead_value_26;
  wire                _zz_io_swRead_value_27;
  wire       [19:0]   _zz_io_swRead_value_28;
  wire       [19:0]   _zz_io_swRead_value_29;
  wire       [19:0]   _zz_io_swRead_value_30;
  wire       [19:0]   _zz_io_swRead_value_31;
  wire                _zz_io_swRead_value_32;
  wire                _zz_io_swRead_value_33;
  wire                _zz_io_swRead_value_34;
  wire                _zz_io_swRead_value_35;
  wire                _zz_io_csrWrite_asid_1;
  wire       [3:0]    _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire       [3:0]    _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_when_TLB_l130;
  wire       [3:0]    _zz_11;
  wire                _zz_when_TLB_l130_1;
  wire                _zz_when_TLB_l130_2;
  wire                when_TLB_l130;
  `ifndef SYNTHESIS
  reg [39:0] io_ctrl_op_string;
  `endif

  function  zz_replaceCounter_willIncrement(input dummy);
    begin
      zz_replaceCounter_willIncrement = 1'b0;
      zz_replaceCounter_willIncrement = 1'b1;
    end
  endfunction
  wire  _zz_12;

  assign _zz_replaceCounter_valueNext_1 = replaceCounter_willIncrement;
  assign _zz_replaceCounter_valueNext = {1'd0, _zz_replaceCounter_valueNext_1};
  assign _zz__zz_when_TLB_l130_2_1 = ((_zz__zz_when_TLB_l130_2_2 == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz__zz_io_csrWrite_asid_1_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_4_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_8_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_9_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_10_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_11_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_12_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_13_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_15_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_17_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_18_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_19_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_20_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_21_1 = _zz_io_csrWrite_asid;
  assign _zz__zz_io_swRead_value_23_1 = _zz_io_csrWrite_asid;
  always @(*) begin
    case(_zz_io_iCacheReq_pageInfo_ppn_4)
      2'b00 : begin
        _zz__zz_io_iCacheReq_pageInfo_ppn_5 = _zz_io_iCacheReq_hit_3;
        _zz__zz_io_iCacheReq_pageInfo_ppn_6 = ((tlbStorage_0_ps == 6'h0c) ? io_iCacheReq_virtPageNumber[0] : io_iCacheReq_virtPageNumber[9]);
        _zz_io_iCacheReq_pageInfo_ppn_7 = tlbStorage_0_pp1_ppn;
        _zz_io_iCacheReq_pageInfo_ppn_8 = tlbStorage_0_pp0_ppn;
        _zz_io_iCacheReq_pageInfo_plv_1 = tlbStorage_0_pp1_plv;
        _zz_io_iCacheReq_pageInfo_plv_2 = tlbStorage_0_pp0_plv;
        _zz_io_iCacheReq_pageInfo_mat_3 = tlbStorage_0_pp1_mat;
        _zz_io_iCacheReq_pageInfo_mat_4 = tlbStorage_0_pp0_mat;
        _zz_io_iCacheReq_pageInfo_d = tlbStorage_0_pp1_d;
        _zz_io_iCacheReq_pageInfo_d_1 = tlbStorage_0_pp0_d;
        _zz_io_iCacheReq_pageInfo_v = tlbStorage_0_pp1_v;
        _zz_io_iCacheReq_pageInfo_v_1 = tlbStorage_0_pp0_v;
      end
      2'b01 : begin
        _zz__zz_io_iCacheReq_pageInfo_ppn_5 = _zz_io_iCacheReq_hit_4;
        _zz__zz_io_iCacheReq_pageInfo_ppn_6 = ((tlbStorage_1_ps == 6'h0c) ? io_iCacheReq_virtPageNumber[0] : io_iCacheReq_virtPageNumber[9]);
        _zz_io_iCacheReq_pageInfo_ppn_7 = tlbStorage_1_pp1_ppn;
        _zz_io_iCacheReq_pageInfo_ppn_8 = tlbStorage_1_pp0_ppn;
        _zz_io_iCacheReq_pageInfo_plv_1 = tlbStorage_1_pp1_plv;
        _zz_io_iCacheReq_pageInfo_plv_2 = tlbStorage_1_pp0_plv;
        _zz_io_iCacheReq_pageInfo_mat_3 = tlbStorage_1_pp1_mat;
        _zz_io_iCacheReq_pageInfo_mat_4 = tlbStorage_1_pp0_mat;
        _zz_io_iCacheReq_pageInfo_d = tlbStorage_1_pp1_d;
        _zz_io_iCacheReq_pageInfo_d_1 = tlbStorage_1_pp0_d;
        _zz_io_iCacheReq_pageInfo_v = tlbStorage_1_pp1_v;
        _zz_io_iCacheReq_pageInfo_v_1 = tlbStorage_1_pp0_v;
      end
      2'b10 : begin
        _zz__zz_io_iCacheReq_pageInfo_ppn_5 = _zz_io_iCacheReq_hit_5;
        _zz__zz_io_iCacheReq_pageInfo_ppn_6 = ((tlbStorage_2_ps == 6'h0c) ? io_iCacheReq_virtPageNumber[0] : io_iCacheReq_virtPageNumber[9]);
        _zz_io_iCacheReq_pageInfo_ppn_7 = tlbStorage_2_pp1_ppn;
        _zz_io_iCacheReq_pageInfo_ppn_8 = tlbStorage_2_pp0_ppn;
        _zz_io_iCacheReq_pageInfo_plv_1 = tlbStorage_2_pp1_plv;
        _zz_io_iCacheReq_pageInfo_plv_2 = tlbStorage_2_pp0_plv;
        _zz_io_iCacheReq_pageInfo_mat_3 = tlbStorage_2_pp1_mat;
        _zz_io_iCacheReq_pageInfo_mat_4 = tlbStorage_2_pp0_mat;
        _zz_io_iCacheReq_pageInfo_d = tlbStorage_2_pp1_d;
        _zz_io_iCacheReq_pageInfo_d_1 = tlbStorage_2_pp0_d;
        _zz_io_iCacheReq_pageInfo_v = tlbStorage_2_pp1_v;
        _zz_io_iCacheReq_pageInfo_v_1 = tlbStorage_2_pp0_v;
      end
      default : begin
        _zz__zz_io_iCacheReq_pageInfo_ppn_5 = _zz_io_iCacheReq_hit_6;
        _zz__zz_io_iCacheReq_pageInfo_ppn_6 = ((tlbStorage_3_ps == 6'h0c) ? io_iCacheReq_virtPageNumber[0] : io_iCacheReq_virtPageNumber[9]);
        _zz_io_iCacheReq_pageInfo_ppn_7 = tlbStorage_3_pp1_ppn;
        _zz_io_iCacheReq_pageInfo_ppn_8 = tlbStorage_3_pp0_ppn;
        _zz_io_iCacheReq_pageInfo_plv_1 = tlbStorage_3_pp1_plv;
        _zz_io_iCacheReq_pageInfo_plv_2 = tlbStorage_3_pp0_plv;
        _zz_io_iCacheReq_pageInfo_mat_3 = tlbStorage_3_pp1_mat;
        _zz_io_iCacheReq_pageInfo_mat_4 = tlbStorage_3_pp0_mat;
        _zz_io_iCacheReq_pageInfo_d = tlbStorage_3_pp1_d;
        _zz_io_iCacheReq_pageInfo_d_1 = tlbStorage_3_pp0_d;
        _zz_io_iCacheReq_pageInfo_v = tlbStorage_3_pp1_v;
        _zz_io_iCacheReq_pageInfo_v_1 = tlbStorage_3_pp0_v;
      end
    endcase
  end

  always @(*) begin
    case(_zz_io_dCacheReq_pageInfo_ppn_2)
      2'b00 : begin
        _zz__zz_io_dCacheReq_pageInfo_ppn_3 = _zz_io_dCacheReq_hit_3;
        _zz__zz_io_dCacheReq_pageInfo_ppn_4 = ((tlbStorage_0_ps == 6'h0c) ? io_dCacheReq_virtPageNumber[0] : io_dCacheReq_virtPageNumber[9]);
        _zz_io_dCacheReq_pageInfo_ppn_5 = tlbStorage_0_pp1_ppn;
        _zz_io_dCacheReq_pageInfo_ppn_6 = tlbStorage_0_pp0_ppn;
        _zz_io_dCacheReq_pageInfo_plv = tlbStorage_0_pp1_plv;
        _zz_io_dCacheReq_pageInfo_plv_1 = tlbStorage_0_pp0_plv;
        _zz_io_dCacheReq_pageInfo_mat_1 = tlbStorage_0_pp1_mat;
        _zz_io_dCacheReq_pageInfo_mat_2 = tlbStorage_0_pp0_mat;
        _zz_io_dCacheReq_pageInfo_d = tlbStorage_0_pp1_d;
        _zz_io_dCacheReq_pageInfo_d_1 = tlbStorage_0_pp0_d;
        _zz_io_dCacheReq_pageInfo_v = tlbStorage_0_pp1_v;
        _zz_io_dCacheReq_pageInfo_v_1 = tlbStorage_0_pp0_v;
      end
      2'b01 : begin
        _zz__zz_io_dCacheReq_pageInfo_ppn_3 = _zz_io_dCacheReq_hit_4;
        _zz__zz_io_dCacheReq_pageInfo_ppn_4 = ((tlbStorage_1_ps == 6'h0c) ? io_dCacheReq_virtPageNumber[0] : io_dCacheReq_virtPageNumber[9]);
        _zz_io_dCacheReq_pageInfo_ppn_5 = tlbStorage_1_pp1_ppn;
        _zz_io_dCacheReq_pageInfo_ppn_6 = tlbStorage_1_pp0_ppn;
        _zz_io_dCacheReq_pageInfo_plv = tlbStorage_1_pp1_plv;
        _zz_io_dCacheReq_pageInfo_plv_1 = tlbStorage_1_pp0_plv;
        _zz_io_dCacheReq_pageInfo_mat_1 = tlbStorage_1_pp1_mat;
        _zz_io_dCacheReq_pageInfo_mat_2 = tlbStorage_1_pp0_mat;
        _zz_io_dCacheReq_pageInfo_d = tlbStorage_1_pp1_d;
        _zz_io_dCacheReq_pageInfo_d_1 = tlbStorage_1_pp0_d;
        _zz_io_dCacheReq_pageInfo_v = tlbStorage_1_pp1_v;
        _zz_io_dCacheReq_pageInfo_v_1 = tlbStorage_1_pp0_v;
      end
      2'b10 : begin
        _zz__zz_io_dCacheReq_pageInfo_ppn_3 = _zz_io_dCacheReq_hit_5;
        _zz__zz_io_dCacheReq_pageInfo_ppn_4 = ((tlbStorage_2_ps == 6'h0c) ? io_dCacheReq_virtPageNumber[0] : io_dCacheReq_virtPageNumber[9]);
        _zz_io_dCacheReq_pageInfo_ppn_5 = tlbStorage_2_pp1_ppn;
        _zz_io_dCacheReq_pageInfo_ppn_6 = tlbStorage_2_pp0_ppn;
        _zz_io_dCacheReq_pageInfo_plv = tlbStorage_2_pp1_plv;
        _zz_io_dCacheReq_pageInfo_plv_1 = tlbStorage_2_pp0_plv;
        _zz_io_dCacheReq_pageInfo_mat_1 = tlbStorage_2_pp1_mat;
        _zz_io_dCacheReq_pageInfo_mat_2 = tlbStorage_2_pp0_mat;
        _zz_io_dCacheReq_pageInfo_d = tlbStorage_2_pp1_d;
        _zz_io_dCacheReq_pageInfo_d_1 = tlbStorage_2_pp0_d;
        _zz_io_dCacheReq_pageInfo_v = tlbStorage_2_pp1_v;
        _zz_io_dCacheReq_pageInfo_v_1 = tlbStorage_2_pp0_v;
      end
      default : begin
        _zz__zz_io_dCacheReq_pageInfo_ppn_3 = _zz_io_dCacheReq_hit_6;
        _zz__zz_io_dCacheReq_pageInfo_ppn_4 = ((tlbStorage_3_ps == 6'h0c) ? io_dCacheReq_virtPageNumber[0] : io_dCacheReq_virtPageNumber[9]);
        _zz_io_dCacheReq_pageInfo_ppn_5 = tlbStorage_3_pp1_ppn;
        _zz_io_dCacheReq_pageInfo_ppn_6 = tlbStorage_3_pp0_ppn;
        _zz_io_dCacheReq_pageInfo_plv = tlbStorage_3_pp1_plv;
        _zz_io_dCacheReq_pageInfo_plv_1 = tlbStorage_3_pp0_plv;
        _zz_io_dCacheReq_pageInfo_mat_1 = tlbStorage_3_pp1_mat;
        _zz_io_dCacheReq_pageInfo_mat_2 = tlbStorage_3_pp0_mat;
        _zz_io_dCacheReq_pageInfo_d = tlbStorage_3_pp1_d;
        _zz_io_dCacheReq_pageInfo_d_1 = tlbStorage_3_pp0_d;
        _zz_io_dCacheReq_pageInfo_v = tlbStorage_3_pp1_v;
        _zz_io_dCacheReq_pageInfo_v_1 = tlbStorage_3_pp0_v;
      end
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_csrWrite_asid_1_1)
      2'b00 : _zz__zz_io_csrWrite_asid_1 = tlbStorage_0_e;
      2'b01 : _zz__zz_io_csrWrite_asid_1 = tlbStorage_1_e;
      2'b10 : _zz__zz_io_csrWrite_asid_1 = tlbStorage_2_e;
      default : _zz__zz_io_csrWrite_asid_1 = tlbStorage_3_e;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_4_1)
      2'b00 : _zz__zz_io_swRead_value_4 = tlbStorage_0_ps;
      2'b01 : _zz__zz_io_swRead_value_4 = tlbStorage_1_ps;
      2'b10 : _zz__zz_io_swRead_value_4 = tlbStorage_2_ps;
      default : _zz__zz_io_swRead_value_4 = tlbStorage_3_ps;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_8_1)
      2'b00 : _zz__zz_io_swRead_value_8 = tlbStorage_0_vppn;
      2'b01 : _zz__zz_io_swRead_value_8 = tlbStorage_1_vppn;
      2'b10 : _zz__zz_io_swRead_value_8 = tlbStorage_2_vppn;
      default : _zz__zz_io_swRead_value_8 = tlbStorage_3_vppn;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_9_1)
      2'b00 : _zz__zz_io_swRead_value_9 = tlbStorage_0_pp0_v;
      2'b01 : _zz__zz_io_swRead_value_9 = tlbStorage_1_pp0_v;
      2'b10 : _zz__zz_io_swRead_value_9 = tlbStorage_2_pp0_v;
      default : _zz__zz_io_swRead_value_9 = tlbStorage_3_pp0_v;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_10_1)
      2'b00 : _zz__zz_io_swRead_value_10 = tlbStorage_0_pp0_d;
      2'b01 : _zz__zz_io_swRead_value_10 = tlbStorage_1_pp0_d;
      2'b10 : _zz__zz_io_swRead_value_10 = tlbStorage_2_pp0_d;
      default : _zz__zz_io_swRead_value_10 = tlbStorage_3_pp0_d;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_11_1)
      2'b00 : _zz__zz_io_swRead_value_11 = tlbStorage_0_pp0_plv;
      2'b01 : _zz__zz_io_swRead_value_11 = tlbStorage_1_pp0_plv;
      2'b10 : _zz__zz_io_swRead_value_11 = tlbStorage_2_pp0_plv;
      default : _zz__zz_io_swRead_value_11 = tlbStorage_3_pp0_plv;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_12_1)
      2'b00 : _zz__zz_io_swRead_value_12 = tlbStorage_0_pp0_mat;
      2'b01 : _zz__zz_io_swRead_value_12 = tlbStorage_1_pp0_mat;
      2'b10 : _zz__zz_io_swRead_value_12 = tlbStorage_2_pp0_mat;
      default : _zz__zz_io_swRead_value_12 = tlbStorage_3_pp0_mat;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_13_1)
      2'b00 : _zz__zz_io_swRead_value_13 = tlbStorage_0_g;
      2'b01 : _zz__zz_io_swRead_value_13 = tlbStorage_1_g;
      2'b10 : _zz__zz_io_swRead_value_13 = tlbStorage_2_g;
      default : _zz__zz_io_swRead_value_13 = tlbStorage_3_g;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_15_1)
      2'b00 : _zz__zz_io_swRead_value_15 = tlbStorage_0_pp0_ppn;
      2'b01 : _zz__zz_io_swRead_value_15 = tlbStorage_1_pp0_ppn;
      2'b10 : _zz__zz_io_swRead_value_15 = tlbStorage_2_pp0_ppn;
      default : _zz__zz_io_swRead_value_15 = tlbStorage_3_pp0_ppn;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_17_1)
      2'b00 : _zz__zz_io_swRead_value_17 = tlbStorage_0_pp1_v;
      2'b01 : _zz__zz_io_swRead_value_17 = tlbStorage_1_pp1_v;
      2'b10 : _zz__zz_io_swRead_value_17 = tlbStorage_2_pp1_v;
      default : _zz__zz_io_swRead_value_17 = tlbStorage_3_pp1_v;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_18_1)
      2'b00 : _zz__zz_io_swRead_value_18 = tlbStorage_0_pp1_d;
      2'b01 : _zz__zz_io_swRead_value_18 = tlbStorage_1_pp1_d;
      2'b10 : _zz__zz_io_swRead_value_18 = tlbStorage_2_pp1_d;
      default : _zz__zz_io_swRead_value_18 = tlbStorage_3_pp1_d;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_19_1)
      2'b00 : _zz__zz_io_swRead_value_19 = tlbStorage_0_pp1_plv;
      2'b01 : _zz__zz_io_swRead_value_19 = tlbStorage_1_pp1_plv;
      2'b10 : _zz__zz_io_swRead_value_19 = tlbStorage_2_pp1_plv;
      default : _zz__zz_io_swRead_value_19 = tlbStorage_3_pp1_plv;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_20_1)
      2'b00 : _zz__zz_io_swRead_value_20 = tlbStorage_0_pp1_mat;
      2'b01 : _zz__zz_io_swRead_value_20 = tlbStorage_1_pp1_mat;
      2'b10 : _zz__zz_io_swRead_value_20 = tlbStorage_2_pp1_mat;
      default : _zz__zz_io_swRead_value_20 = tlbStorage_3_pp1_mat;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_21_1)
      2'b00 : _zz__zz_io_swRead_value_21 = tlbStorage_0_g;
      2'b01 : _zz__zz_io_swRead_value_21 = tlbStorage_1_g;
      2'b10 : _zz__zz_io_swRead_value_21 = tlbStorage_2_g;
      default : _zz__zz_io_swRead_value_21 = tlbStorage_3_g;
    endcase
  end

  always @(*) begin
    case(_zz__zz_io_swRead_value_23_1)
      2'b00 : _zz__zz_io_swRead_value_23 = tlbStorage_0_pp1_ppn;
      2'b01 : _zz__zz_io_swRead_value_23 = tlbStorage_1_pp1_ppn;
      2'b10 : _zz__zz_io_swRead_value_23 = tlbStorage_2_pp1_ppn;
      default : _zz__zz_io_swRead_value_23 = tlbStorage_3_pp1_ppn;
    endcase
  end

  always @(*) begin
    case(io_ctrl_index)
      2'b00 : begin
        _zz__zz_when_TLB_l130 = tlbStorage_0_g;
        _zz__zz_when_TLB_l130_1 = tlbStorage_0_asid;
        _zz__zz_when_TLB_l130_2 = tlbStorage_0_vppn;
        _zz__zz_when_TLB_l130_2_2 = tlbStorage_0_ps;
      end
      2'b01 : begin
        _zz__zz_when_TLB_l130 = tlbStorage_1_g;
        _zz__zz_when_TLB_l130_1 = tlbStorage_1_asid;
        _zz__zz_when_TLB_l130_2 = tlbStorage_1_vppn;
        _zz__zz_when_TLB_l130_2_2 = tlbStorage_1_ps;
      end
      2'b10 : begin
        _zz__zz_when_TLB_l130 = tlbStorage_2_g;
        _zz__zz_when_TLB_l130_1 = tlbStorage_2_asid;
        _zz__zz_when_TLB_l130_2 = tlbStorage_2_vppn;
        _zz__zz_when_TLB_l130_2_2 = tlbStorage_2_ps;
      end
      default : begin
        _zz__zz_when_TLB_l130 = tlbStorage_3_g;
        _zz__zz_when_TLB_l130_1 = tlbStorage_3_asid;
        _zz__zz_when_TLB_l130_2 = tlbStorage_3_vppn;
        _zz__zz_when_TLB_l130_2_2 = tlbStorage_3_ps;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_ctrl_op)
      TLBOp_nop : io_ctrl_op_string = "nop  ";
      TLBOp_srch : io_ctrl_op_string = "srch ";
      TLBOp_read : io_ctrl_op_string = "read ";
      TLBOp_write : io_ctrl_op_string = "write";
      TLBOp_fill : io_ctrl_op_string = "fill ";
      TLBOp_inv : io_ctrl_op_string = "inv  ";
      default : io_ctrl_op_string = "?????";
    endcase
  end
  `endif

  assign when_TLB_l177 = (_zz_when_TLB_l177_1 && (! _zz_when_TLB_l177));
  assign when_TLB_l178 = ((io_iCacheReq_virtPageNumber[19 : 17] == _zz_when_TLB_l178_2) && (((_zz_io_iCacheReq_pageInfo_plv == 2'b11) && _zz_when_TLB_l178_1) || ((_zz_io_iCacheReq_pageInfo_plv == 2'b00) && _zz_when_TLB_l178)));
  always @(*) begin
    if(when_TLB_l177) begin
      if(when_TLB_l178) begin
        io_iCacheReq_pageInfo_ppn = {_zz_io_iCacheReq_pageInfo_ppn,io_iCacheReq_virtPageNumber[16 : 0]};
      end else begin
        if(when_TLB_l185) begin
          io_iCacheReq_pageInfo_ppn = {_zz_io_iCacheReq_pageInfo_ppn_1,io_iCacheReq_virtPageNumber[16 : 0]};
        end else begin
          io_iCacheReq_pageInfo_ppn = (((_zz_io_iCacheReq_pageInfo_ppn_6 ? _zz_io_iCacheReq_pageInfo_ppn_7 : _zz_io_iCacheReq_pageInfo_ppn_8) & (~ _zz_io_iCacheReq_pageInfo_ppn_5)) | (io_iCacheReq_virtPageNumber & _zz_io_iCacheReq_pageInfo_ppn_5));
        end
      end
    end else begin
      if(when_TLB_l195) begin
        io_iCacheReq_pageInfo_ppn = io_iCacheReq_virtPageNumber;
      end else begin
        io_iCacheReq_pageInfo_ppn = io_iCacheReq_virtPageNumber;
      end
    end
  end

  always @(*) begin
    if(when_TLB_l177) begin
      if(when_TLB_l178) begin
        io_iCacheReq_pageInfo_plv = _zz_io_iCacheReq_pageInfo_plv;
      end else begin
        if(when_TLB_l185) begin
          io_iCacheReq_pageInfo_plv = _zz_io_iCacheReq_pageInfo_plv;
        end else begin
          io_iCacheReq_pageInfo_plv = (_zz_io_iCacheReq_pageInfo_ppn_6 ? _zz_io_iCacheReq_pageInfo_plv_1 : _zz_io_iCacheReq_pageInfo_plv_2);
        end
      end
    end else begin
      if(when_TLB_l195) begin
        io_iCacheReq_pageInfo_plv = _zz_io_iCacheReq_pageInfo_plv;
      end else begin
        io_iCacheReq_pageInfo_plv = _zz_io_iCacheReq_pageInfo_plv;
      end
    end
  end

  always @(*) begin
    if(when_TLB_l177) begin
      if(when_TLB_l178) begin
        io_iCacheReq_pageInfo_mat = _zz_io_iCacheReq_pageInfo_mat_1;
      end else begin
        if(when_TLB_l185) begin
          io_iCacheReq_pageInfo_mat = _zz_io_iCacheReq_pageInfo_mat_2;
        end else begin
          io_iCacheReq_pageInfo_mat = (_zz_io_iCacheReq_pageInfo_ppn_6 ? _zz_io_iCacheReq_pageInfo_mat_3 : _zz_io_iCacheReq_pageInfo_mat_4);
        end
      end
    end else begin
      if(when_TLB_l195) begin
        io_iCacheReq_pageInfo_mat = _zz_io_iCacheReq_pageInfo_mat;
      end else begin
        io_iCacheReq_pageInfo_mat = _zz_io_iCacheReq_pageInfo_mat;
      end
    end
  end

  always @(*) begin
    if(when_TLB_l177) begin
      if(when_TLB_l178) begin
        io_iCacheReq_pageInfo_d = 1'b1;
      end else begin
        if(when_TLB_l185) begin
          io_iCacheReq_pageInfo_d = 1'b1;
        end else begin
          io_iCacheReq_pageInfo_d = (_zz_io_iCacheReq_pageInfo_ppn_6 ? _zz_io_iCacheReq_pageInfo_d : _zz_io_iCacheReq_pageInfo_d_1);
        end
      end
    end else begin
      if(when_TLB_l195) begin
        io_iCacheReq_pageInfo_d = 1'b1;
      end else begin
        io_iCacheReq_pageInfo_d = 1'b1;
      end
    end
  end

  always @(*) begin
    if(when_TLB_l177) begin
      if(when_TLB_l178) begin
        io_iCacheReq_pageInfo_v = 1'b1;
      end else begin
        if(when_TLB_l185) begin
          io_iCacheReq_pageInfo_v = 1'b1;
        end else begin
          io_iCacheReq_pageInfo_v = (_zz_io_iCacheReq_pageInfo_ppn_6 ? _zz_io_iCacheReq_pageInfo_v : _zz_io_iCacheReq_pageInfo_v_1);
        end
      end
    end else begin
      if(when_TLB_l195) begin
        io_iCacheReq_pageInfo_v = 1'b1;
      end else begin
        io_iCacheReq_pageInfo_v = 1'b1;
      end
    end
  end

  always @(*) begin
    if(when_TLB_l177) begin
      if(when_TLB_l178) begin
        io_iCacheReq_hit = 1'b1;
      end else begin
        if(when_TLB_l185) begin
          io_iCacheReq_hit = 1'b1;
        end else begin
          io_iCacheReq_hit = ((((1'b0 || ((((tlbStorage_0_g || (tlbStorage_0_asid == io_csrInfo_asid)) && tlbStorage_0_e) && ((tlbStorage_0_vppn ^ _zz_io_iCacheReq_hit_3[19 : 1]) == (io_iCacheReq_virtPageNumber[19 : 1] ^ _zz_io_iCacheReq_hit_3[19 : 1]))) == _zz_io_iCacheReq_hit_7)) || (_zz_io_iCacheReq_hit == _zz_io_iCacheReq_hit_7)) || (_zz_io_iCacheReq_hit_1 == _zz_io_iCacheReq_hit_7)) || (_zz_io_iCacheReq_hit_2 == _zz_io_iCacheReq_hit_7));
        end
      end
    end else begin
      if(when_TLB_l195) begin
        io_iCacheReq_hit = 1'b1;
      end else begin
        io_iCacheReq_hit = 1'b1;
      end
    end
  end

  assign _zz_io_iCacheReq_hit_3 = ((tlbStorage_0_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_iCacheReq_hit = (((tlbStorage_1_g || (tlbStorage_1_asid == io_csrInfo_asid)) && tlbStorage_1_e) && ((tlbStorage_1_vppn ^ _zz_io_iCacheReq_hit_4[19 : 1]) == (io_iCacheReq_virtPageNumber[19 : 1] ^ _zz_io_iCacheReq_hit_4[19 : 1])));
  assign _zz_io_iCacheReq_hit_4 = ((tlbStorage_1_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_iCacheReq_hit_1 = (((tlbStorage_2_g || (tlbStorage_2_asid == io_csrInfo_asid)) && tlbStorage_2_e) && ((tlbStorage_2_vppn ^ _zz_io_iCacheReq_hit_5[19 : 1]) == (io_iCacheReq_virtPageNumber[19 : 1] ^ _zz_io_iCacheReq_hit_5[19 : 1])));
  assign _zz_io_iCacheReq_hit_5 = ((tlbStorage_2_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_iCacheReq_hit_2 = (((tlbStorage_3_g || (tlbStorage_3_asid == io_csrInfo_asid)) && tlbStorage_3_e) && ((tlbStorage_3_vppn ^ _zz_io_iCacheReq_hit_6[19 : 1]) == (io_iCacheReq_virtPageNumber[19 : 1] ^ _zz_io_iCacheReq_hit_6[19 : 1])));
  assign _zz_io_iCacheReq_hit_6 = ((tlbStorage_3_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_iCacheReq_pageInfo_ppn_2 = (_zz_io_iCacheReq_hit || _zz_io_iCacheReq_hit_2);
  assign _zz_io_iCacheReq_pageInfo_ppn_3 = (_zz_io_iCacheReq_hit_1 || _zz_io_iCacheReq_hit_2);
  assign _zz_io_iCacheReq_pageInfo_ppn_4 = {_zz_io_iCacheReq_pageInfo_ppn_3,_zz_io_iCacheReq_pageInfo_ppn_2};
  assign _zz_io_iCacheReq_pageInfo_ppn_5 = _zz__zz_io_iCacheReq_pageInfo_ppn_5;
  assign _zz_io_iCacheReq_pageInfo_ppn_6 = _zz__zz_io_iCacheReq_pageInfo_ppn_6;
  assign _zz_io_iCacheReq_hit_7 = 1'b1;
  assign when_TLB_l185 = ((io_iCacheReq_virtPageNumber[19 : 17] == _zz_when_TLB_l185_2) && (((_zz_io_iCacheReq_pageInfo_plv == 2'b11) && _zz_when_TLB_l185_1) || ((_zz_io_iCacheReq_pageInfo_plv == 2'b00) && _zz_when_TLB_l185)));
  assign when_TLB_l195 = ((! _zz_when_TLB_l177_1) && _zz_when_TLB_l177);
  assign when_TLB_l177_1 = (_zz_when_TLB_l177_1 && (! _zz_when_TLB_l177));
  assign when_TLB_l178_1 = ((io_dCacheReq_virtPageNumber[19 : 17] == _zz_when_TLB_l178_2) && (((_zz_io_iCacheReq_pageInfo_plv == 2'b11) && _zz_when_TLB_l178_1) || ((_zz_io_iCacheReq_pageInfo_plv == 2'b00) && _zz_when_TLB_l178)));
  always @(*) begin
    if(when_TLB_l177_1) begin
      if(when_TLB_l178_1) begin
        io_dCacheReq_pageInfo_ppn = {_zz_io_iCacheReq_pageInfo_ppn,io_dCacheReq_virtPageNumber[16 : 0]};
      end else begin
        if(when_TLB_l185_1) begin
          io_dCacheReq_pageInfo_ppn = {_zz_io_iCacheReq_pageInfo_ppn_1,io_dCacheReq_virtPageNumber[16 : 0]};
        end else begin
          io_dCacheReq_pageInfo_ppn = (((_zz_io_dCacheReq_pageInfo_ppn_4 ? _zz_io_dCacheReq_pageInfo_ppn_5 : _zz_io_dCacheReq_pageInfo_ppn_6) & (~ _zz_io_dCacheReq_pageInfo_ppn_3)) | (io_dCacheReq_virtPageNumber & _zz_io_dCacheReq_pageInfo_ppn_3));
        end
      end
    end else begin
      if(when_TLB_l195_1) begin
        io_dCacheReq_pageInfo_ppn = io_dCacheReq_virtPageNumber;
      end else begin
        io_dCacheReq_pageInfo_ppn = io_dCacheReq_virtPageNumber;
      end
    end
  end

  always @(*) begin
    if(when_TLB_l177_1) begin
      if(when_TLB_l178_1) begin
        io_dCacheReq_pageInfo_plv = _zz_io_iCacheReq_pageInfo_plv;
      end else begin
        if(when_TLB_l185_1) begin
          io_dCacheReq_pageInfo_plv = _zz_io_iCacheReq_pageInfo_plv;
        end else begin
          io_dCacheReq_pageInfo_plv = (_zz_io_dCacheReq_pageInfo_ppn_4 ? _zz_io_dCacheReq_pageInfo_plv : _zz_io_dCacheReq_pageInfo_plv_1);
        end
      end
    end else begin
      if(when_TLB_l195_1) begin
        io_dCacheReq_pageInfo_plv = _zz_io_iCacheReq_pageInfo_plv;
      end else begin
        io_dCacheReq_pageInfo_plv = _zz_io_iCacheReq_pageInfo_plv;
      end
    end
  end

  always @(*) begin
    if(when_TLB_l177_1) begin
      if(when_TLB_l178_1) begin
        io_dCacheReq_pageInfo_mat = _zz_io_iCacheReq_pageInfo_mat_1;
      end else begin
        if(when_TLB_l185_1) begin
          io_dCacheReq_pageInfo_mat = _zz_io_iCacheReq_pageInfo_mat_2;
        end else begin
          io_dCacheReq_pageInfo_mat = (_zz_io_dCacheReq_pageInfo_ppn_4 ? _zz_io_dCacheReq_pageInfo_mat_1 : _zz_io_dCacheReq_pageInfo_mat_2);
        end
      end
    end else begin
      if(when_TLB_l195_1) begin
        io_dCacheReq_pageInfo_mat = _zz_io_dCacheReq_pageInfo_mat;
      end else begin
        io_dCacheReq_pageInfo_mat = _zz_io_dCacheReq_pageInfo_mat;
      end
    end
  end

  always @(*) begin
    if(when_TLB_l177_1) begin
      if(when_TLB_l178_1) begin
        io_dCacheReq_pageInfo_d = 1'b1;
      end else begin
        if(when_TLB_l185_1) begin
          io_dCacheReq_pageInfo_d = 1'b1;
        end else begin
          io_dCacheReq_pageInfo_d = (_zz_io_dCacheReq_pageInfo_ppn_4 ? _zz_io_dCacheReq_pageInfo_d : _zz_io_dCacheReq_pageInfo_d_1);
        end
      end
    end else begin
      if(when_TLB_l195_1) begin
        io_dCacheReq_pageInfo_d = 1'b1;
      end else begin
        io_dCacheReq_pageInfo_d = 1'b1;
      end
    end
  end

  always @(*) begin
    if(when_TLB_l177_1) begin
      if(when_TLB_l178_1) begin
        io_dCacheReq_pageInfo_v = 1'b1;
      end else begin
        if(when_TLB_l185_1) begin
          io_dCacheReq_pageInfo_v = 1'b1;
        end else begin
          io_dCacheReq_pageInfo_v = (_zz_io_dCacheReq_pageInfo_ppn_4 ? _zz_io_dCacheReq_pageInfo_v : _zz_io_dCacheReq_pageInfo_v_1);
        end
      end
    end else begin
      if(when_TLB_l195_1) begin
        io_dCacheReq_pageInfo_v = 1'b1;
      end else begin
        io_dCacheReq_pageInfo_v = 1'b1;
      end
    end
  end

  always @(*) begin
    if(when_TLB_l177_1) begin
      if(when_TLB_l178_1) begin
        io_dCacheReq_hit = 1'b1;
      end else begin
        if(when_TLB_l185_1) begin
          io_dCacheReq_hit = 1'b1;
        end else begin
          io_dCacheReq_hit = ((((1'b0 || ((((tlbStorage_0_g || (tlbStorage_0_asid == io_csrInfo_asid)) && tlbStorage_0_e) && ((tlbStorage_0_vppn ^ _zz_io_dCacheReq_hit_3[19 : 1]) == (io_dCacheReq_virtPageNumber[19 : 1] ^ _zz_io_dCacheReq_hit_3[19 : 1]))) == _zz_io_dCacheReq_hit_7)) || (_zz_io_dCacheReq_hit == _zz_io_dCacheReq_hit_7)) || (_zz_io_dCacheReq_hit_1 == _zz_io_dCacheReq_hit_7)) || (_zz_io_dCacheReq_hit_2 == _zz_io_dCacheReq_hit_7));
        end
      end
    end else begin
      if(when_TLB_l195_1) begin
        io_dCacheReq_hit = 1'b1;
      end else begin
        io_dCacheReq_hit = 1'b1;
      end
    end
  end

  assign _zz_io_dCacheReq_hit_3 = ((tlbStorage_0_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_dCacheReq_hit = (((tlbStorage_1_g || (tlbStorage_1_asid == io_csrInfo_asid)) && tlbStorage_1_e) && ((tlbStorage_1_vppn ^ _zz_io_dCacheReq_hit_4[19 : 1]) == (io_dCacheReq_virtPageNumber[19 : 1] ^ _zz_io_dCacheReq_hit_4[19 : 1])));
  assign _zz_io_dCacheReq_hit_4 = ((tlbStorage_1_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_dCacheReq_hit_1 = (((tlbStorage_2_g || (tlbStorage_2_asid == io_csrInfo_asid)) && tlbStorage_2_e) && ((tlbStorage_2_vppn ^ _zz_io_dCacheReq_hit_5[19 : 1]) == (io_dCacheReq_virtPageNumber[19 : 1] ^ _zz_io_dCacheReq_hit_5[19 : 1])));
  assign _zz_io_dCacheReq_hit_5 = ((tlbStorage_2_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_dCacheReq_hit_2 = (((tlbStorage_3_g || (tlbStorage_3_asid == io_csrInfo_asid)) && tlbStorage_3_e) && ((tlbStorage_3_vppn ^ _zz_io_dCacheReq_hit_6[19 : 1]) == (io_dCacheReq_virtPageNumber[19 : 1] ^ _zz_io_dCacheReq_hit_6[19 : 1])));
  assign _zz_io_dCacheReq_hit_6 = ((tlbStorage_3_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_dCacheReq_pageInfo_ppn = (_zz_io_dCacheReq_hit || _zz_io_dCacheReq_hit_2);
  assign _zz_io_dCacheReq_pageInfo_ppn_1 = (_zz_io_dCacheReq_hit_1 || _zz_io_dCacheReq_hit_2);
  assign _zz_io_dCacheReq_pageInfo_ppn_2 = {_zz_io_dCacheReq_pageInfo_ppn_1,_zz_io_dCacheReq_pageInfo_ppn};
  assign _zz_io_dCacheReq_pageInfo_ppn_3 = _zz__zz_io_dCacheReq_pageInfo_ppn_3;
  assign _zz_io_dCacheReq_pageInfo_ppn_4 = _zz__zz_io_dCacheReq_pageInfo_ppn_4;
  assign _zz_io_dCacheReq_hit_7 = 1'b1;
  assign when_TLB_l185_1 = ((io_dCacheReq_virtPageNumber[19 : 17] == _zz_when_TLB_l185_2) && (((_zz_io_iCacheReq_pageInfo_plv == 2'b11) && _zz_when_TLB_l185_1) || ((_zz_io_iCacheReq_pageInfo_plv == 2'b00) && _zz_when_TLB_l185)));
  assign when_TLB_l195_1 = ((! _zz_when_TLB_l177_1) && _zz_when_TLB_l177);
  always @(*) begin
    io_csrWrite_asid = 10'h000;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        io_csrWrite_asid = (_zz_io_csrWrite_asid_1 ? io_csrInfo_asid : 10'h000);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_2 = 2'b00;
    case(io_ctrl_op)
      TLBOp_srch : begin
        _zz_io_swRead_value_2 = (_zz_io_swRead_value_33 ? {_zz_io_swRead_value_35,_zz_io_swRead_value_34} : _zz_io_csrWrite_asid);
      end
      TLBOp_read : begin
        _zz_io_swRead_value_2 = _zz_io_csrWrite_asid;
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_3 = 22'h000000;
    case(io_ctrl_op)
      TLBOp_srch : begin
        _zz_io_swRead_value_3 = _zz_io_swRead_value;
      end
      TLBOp_read : begin
        _zz_io_swRead_value_3 = _zz_io_swRead_value;
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_4 = 6'h00;
    case(io_ctrl_op)
      TLBOp_srch : begin
        _zz_io_swRead_value_4 = _zz_entryToFill_ps;
      end
      TLBOp_read : begin
        _zz_io_swRead_value_4 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_4 : 6'h00);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_5 = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
        _zz_io_swRead_value_5 = _zz_io_swRead_value_1;
      end
      TLBOp_read : begin
        _zz_io_swRead_value_5 = _zz_io_swRead_value_1;
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_6 = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
        _zz_io_swRead_value_6 = (! _zz_io_swRead_value_33);
      end
      TLBOp_read : begin
        _zz_io_swRead_value_6 = (! _zz_io_csrWrite_asid_1);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_7 = 13'h0000;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_7 = 13'h0000;
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_8 = 19'h00000;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_8 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_8 : 19'h00000);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_9 = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_9 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_9 : 1'b0);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_10 = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_10 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_10 : 1'b0);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_11 = 2'b00;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_11 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_11 : 2'b00);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_12 = 2'b00;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_12 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_12 : 2'b00);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_13 = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_13 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_13 : 1'b0);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_14 = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_14 = 1'b0;
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_15 = 20'h00000;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_15 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_15 : 20'h00000);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_16 = 4'b0000;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_16 = 4'b0000;
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_17 = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_17 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_17 : 1'b0);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_18 = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_18 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_18 : 1'b0);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_19 = 2'b00;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_19 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_19 : 2'b00);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_20 = 2'b00;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_20 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_20 : 2'b00);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_21 = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_21 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_21 : 1'b0);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_22 = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_22 = 1'b0;
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_23 = 20'h00000;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_23 = (_zz_io_csrWrite_asid_1 ? _zz__zz_io_swRead_value_23 : 20'h00000);
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_swRead_value_24 = 4'b0000;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        _zz_io_swRead_value_24 = 4'b0000;
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_csrWrite_idxWen = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
        io_csrWrite_idxWen = 1'b1;
      end
      TLBOp_read : begin
        io_csrWrite_idxWen = 1'b1;
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_csrWrite_entryWen = 1'b0;
    case(io_ctrl_op)
      TLBOp_srch : begin
      end
      TLBOp_read : begin
        io_csrWrite_entryWen = 1'b1;
      end
      TLBOp_write : begin
      end
      TLBOp_fill : begin
      end
      TLBOp_inv : begin
      end
      default : begin
      end
    endcase
  end

  assign entryToFill_vppn = _zz_entryToFill_vppn;
  assign entryToFill_ps = _zz_entryToFill_ps;
  assign entryToFill_g = (_zz_entryToFill_g && _zz_entryToFill_g_1);
  assign entryToFill_asid = io_csrInfo_asid;
  assign entryToFill_e = ((_zz_entryToFill_e == 6'h3f) || (! _zz_entryToFill_e_1));
  assign entryToFill_pp0_ppn = _zz_entryToFill_pp0_ppn;
  assign entryToFill_pp0_plv = _zz_entryToFill_pp0_plv;
  assign entryToFill_pp0_mat = _zz_entryToFill_pp0_mat;
  assign entryToFill_pp0_d = _zz_entryToFill_pp0_d;
  assign entryToFill_pp0_v = _zz_entryToFill_pp0_v;
  assign entryToFill_pp1_ppn = _zz_entryToFill_pp1_ppn;
  assign entryToFill_pp1_plv = _zz_entryToFill_pp1_plv;
  assign entryToFill_pp1_mat = _zz_entryToFill_pp1_mat;
  assign entryToFill_pp1_d = _zz_entryToFill_pp1_d;
  assign entryToFill_pp1_v = _zz_entryToFill_pp1_v;
  assign _zz_12 = zz_replaceCounter_willIncrement(1'b0);
  always @(*) replaceCounter_willIncrement = _zz_12;
  assign replaceCounter_willClear = 1'b0;
  assign replaceCounter_willOverflowIfInc = (replaceCounter_value == 2'b11);
  assign replaceCounter_willOverflow = (replaceCounter_willOverflowIfInc && replaceCounter_willIncrement);
  always @(*) begin
    replaceCounter_valueNext = (replaceCounter_value + _zz_replaceCounter_valueNext);
    if(replaceCounter_willClear) begin
      replaceCounter_valueNext = 2'b00;
    end
  end

  assign _zz_io_swRead_value_32 = 1'b1;
  assign _zz_io_swRead_value_33 = ((((1'b0 || ((((tlbStorage_0_g || (tlbStorage_0_asid == io_csrInfo_asid)) && tlbStorage_0_e) && ((tlbStorage_0_vppn ^ _zz_io_swRead_value_28[19 : 1]) == (_zz_entryToFill_vppn ^ _zz_io_swRead_value_28[19 : 1]))) == _zz_io_swRead_value_32)) || (_zz_io_swRead_value_25 == _zz_io_swRead_value_32)) || (_zz_io_swRead_value_26 == _zz_io_swRead_value_32)) || (_zz_io_swRead_value_27 == _zz_io_swRead_value_32));
  assign _zz_io_swRead_value_28 = ((tlbStorage_0_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_swRead_value_25 = (((tlbStorage_1_g || (tlbStorage_1_asid == io_csrInfo_asid)) && tlbStorage_1_e) && ((tlbStorage_1_vppn ^ _zz_io_swRead_value_29[19 : 1]) == (_zz_entryToFill_vppn ^ _zz_io_swRead_value_29[19 : 1])));
  assign _zz_io_swRead_value_29 = ((tlbStorage_1_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_swRead_value_26 = (((tlbStorage_2_g || (tlbStorage_2_asid == io_csrInfo_asid)) && tlbStorage_2_e) && ((tlbStorage_2_vppn ^ _zz_io_swRead_value_30[19 : 1]) == (_zz_entryToFill_vppn ^ _zz_io_swRead_value_30[19 : 1])));
  assign _zz_io_swRead_value_30 = ((tlbStorage_2_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_swRead_value_27 = (((tlbStorage_3_g || (tlbStorage_3_asid == io_csrInfo_asid)) && tlbStorage_3_e) && ((tlbStorage_3_vppn ^ _zz_io_swRead_value_31[19 : 1]) == (_zz_entryToFill_vppn ^ _zz_io_swRead_value_31[19 : 1])));
  assign _zz_io_swRead_value_31 = ((tlbStorage_3_ps == 6'h0c) ? 20'h00000 : 20'h001ff);
  assign _zz_io_swRead_value_34 = (_zz_io_swRead_value_25 || _zz_io_swRead_value_27);
  assign _zz_io_swRead_value_35 = (_zz_io_swRead_value_26 || _zz_io_swRead_value_27);
  assign _zz_io_csrWrite_asid_1 = _zz__zz_io_csrWrite_asid_1;
  assign _zz_1 = ({3'd0,1'b1} <<< _zz_io_csrWrite_asid);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = ({3'd0,1'b1} <<< replaceCounter_value);
  assign _zz_7 = _zz_6[0];
  assign _zz_8 = _zz_6[1];
  assign _zz_9 = _zz_6[2];
  assign _zz_10 = _zz_6[3];
  assign _zz_when_TLB_l130 = _zz__zz_when_TLB_l130;
  assign _zz_11 = ({3'd0,1'b1} <<< io_ctrl_index);
  assign _zz_when_TLB_l130_1 = (_zz__zz_when_TLB_l130_1 == io_ctrl_asid);
  assign _zz_when_TLB_l130_2 = ((_zz__zz_when_TLB_l130_2 ^ io_ctrl_invVA) == (io_ctrl_invVA ^ _zz__zz_when_TLB_l130_2_1[19 : 1]));
  assign when_TLB_l130 = ((((io_ctrl_invGlobal && _zz_when_TLB_l130) || (io_ctrl_invLocalVAMatch && (((! _zz_when_TLB_l130) && _zz_when_TLB_l130_2) && _zz_when_TLB_l130_1))) || (io_ctrl_invLocalVANotMatch && (((! _zz_when_TLB_l130) && (! _zz_when_TLB_l130_2)) && _zz_when_TLB_l130_1))) || (io_ctrl_invLocal && (! _zz_when_TLB_l130)));
  always @(posedge aclk) begin
    if(!aresetn) begin
      tlbStorage_0_vppn <= 19'h00000;
      tlbStorage_0_ps <= 6'h00;
      tlbStorage_0_g <= 1'b0;
      tlbStorage_0_asid <= 10'h000;
      tlbStorage_0_e <= 1'b0;
      tlbStorage_0_pp0_ppn <= 20'h00000;
      tlbStorage_0_pp0_plv <= 2'b00;
      tlbStorage_0_pp0_mat <= 2'b00;
      tlbStorage_0_pp0_d <= 1'b0;
      tlbStorage_0_pp0_v <= 1'b0;
      tlbStorage_0_pp1_ppn <= 20'h00000;
      tlbStorage_0_pp1_plv <= 2'b00;
      tlbStorage_0_pp1_mat <= 2'b00;
      tlbStorage_0_pp1_d <= 1'b0;
      tlbStorage_0_pp1_v <= 1'b0;
      tlbStorage_1_vppn <= 19'h00000;
      tlbStorage_1_ps <= 6'h00;
      tlbStorage_1_g <= 1'b0;
      tlbStorage_1_asid <= 10'h000;
      tlbStorage_1_e <= 1'b0;
      tlbStorage_1_pp0_ppn <= 20'h00000;
      tlbStorage_1_pp0_plv <= 2'b00;
      tlbStorage_1_pp0_mat <= 2'b00;
      tlbStorage_1_pp0_d <= 1'b0;
      tlbStorage_1_pp0_v <= 1'b0;
      tlbStorage_1_pp1_ppn <= 20'h00000;
      tlbStorage_1_pp1_plv <= 2'b00;
      tlbStorage_1_pp1_mat <= 2'b00;
      tlbStorage_1_pp1_d <= 1'b0;
      tlbStorage_1_pp1_v <= 1'b0;
      tlbStorage_2_vppn <= 19'h00000;
      tlbStorage_2_ps <= 6'h00;
      tlbStorage_2_g <= 1'b0;
      tlbStorage_2_asid <= 10'h000;
      tlbStorage_2_e <= 1'b0;
      tlbStorage_2_pp0_ppn <= 20'h00000;
      tlbStorage_2_pp0_plv <= 2'b00;
      tlbStorage_2_pp0_mat <= 2'b00;
      tlbStorage_2_pp0_d <= 1'b0;
      tlbStorage_2_pp0_v <= 1'b0;
      tlbStorage_2_pp1_ppn <= 20'h00000;
      tlbStorage_2_pp1_plv <= 2'b00;
      tlbStorage_2_pp1_mat <= 2'b00;
      tlbStorage_2_pp1_d <= 1'b0;
      tlbStorage_2_pp1_v <= 1'b0;
      tlbStorage_3_vppn <= 19'h00000;
      tlbStorage_3_ps <= 6'h00;
      tlbStorage_3_g <= 1'b0;
      tlbStorage_3_asid <= 10'h000;
      tlbStorage_3_e <= 1'b0;
      tlbStorage_3_pp0_ppn <= 20'h00000;
      tlbStorage_3_pp0_plv <= 2'b00;
      tlbStorage_3_pp0_mat <= 2'b00;
      tlbStorage_3_pp0_d <= 1'b0;
      tlbStorage_3_pp0_v <= 1'b0;
      tlbStorage_3_pp1_ppn <= 20'h00000;
      tlbStorage_3_pp1_plv <= 2'b00;
      tlbStorage_3_pp1_mat <= 2'b00;
      tlbStorage_3_pp1_d <= 1'b0;
      tlbStorage_3_pp1_v <= 1'b0;
      replaceCounter_value <= 2'b00;
    end else begin
      replaceCounter_value <= replaceCounter_valueNext;
      case(io_ctrl_op)
        TLBOp_srch : begin
        end
        TLBOp_read : begin
        end
        TLBOp_write : begin
          if(_zz_2) begin
            tlbStorage_0_vppn <= entryToFill_vppn;
          end
          if(_zz_3) begin
            tlbStorage_1_vppn <= entryToFill_vppn;
          end
          if(_zz_4) begin
            tlbStorage_2_vppn <= entryToFill_vppn;
          end
          if(_zz_5) begin
            tlbStorage_3_vppn <= entryToFill_vppn;
          end
          if(_zz_2) begin
            tlbStorage_0_ps <= entryToFill_ps;
          end
          if(_zz_3) begin
            tlbStorage_1_ps <= entryToFill_ps;
          end
          if(_zz_4) begin
            tlbStorage_2_ps <= entryToFill_ps;
          end
          if(_zz_5) begin
            tlbStorage_3_ps <= entryToFill_ps;
          end
          if(_zz_2) begin
            tlbStorage_0_g <= entryToFill_g;
          end
          if(_zz_3) begin
            tlbStorage_1_g <= entryToFill_g;
          end
          if(_zz_4) begin
            tlbStorage_2_g <= entryToFill_g;
          end
          if(_zz_5) begin
            tlbStorage_3_g <= entryToFill_g;
          end
          if(_zz_2) begin
            tlbStorage_0_asid <= entryToFill_asid;
          end
          if(_zz_3) begin
            tlbStorage_1_asid <= entryToFill_asid;
          end
          if(_zz_4) begin
            tlbStorage_2_asid <= entryToFill_asid;
          end
          if(_zz_5) begin
            tlbStorage_3_asid <= entryToFill_asid;
          end
          if(_zz_2) begin
            tlbStorage_0_e <= entryToFill_e;
          end
          if(_zz_3) begin
            tlbStorage_1_e <= entryToFill_e;
          end
          if(_zz_4) begin
            tlbStorage_2_e <= entryToFill_e;
          end
          if(_zz_5) begin
            tlbStorage_3_e <= entryToFill_e;
          end
          if(_zz_2) begin
            tlbStorage_0_pp0_ppn <= entryToFill_pp0_ppn;
          end
          if(_zz_3) begin
            tlbStorage_1_pp0_ppn <= entryToFill_pp0_ppn;
          end
          if(_zz_4) begin
            tlbStorage_2_pp0_ppn <= entryToFill_pp0_ppn;
          end
          if(_zz_5) begin
            tlbStorage_3_pp0_ppn <= entryToFill_pp0_ppn;
          end
          if(_zz_2) begin
            tlbStorage_0_pp0_plv <= entryToFill_pp0_plv;
          end
          if(_zz_3) begin
            tlbStorage_1_pp0_plv <= entryToFill_pp0_plv;
          end
          if(_zz_4) begin
            tlbStorage_2_pp0_plv <= entryToFill_pp0_plv;
          end
          if(_zz_5) begin
            tlbStorage_3_pp0_plv <= entryToFill_pp0_plv;
          end
          if(_zz_2) begin
            tlbStorage_0_pp0_mat <= entryToFill_pp0_mat;
          end
          if(_zz_3) begin
            tlbStorage_1_pp0_mat <= entryToFill_pp0_mat;
          end
          if(_zz_4) begin
            tlbStorage_2_pp0_mat <= entryToFill_pp0_mat;
          end
          if(_zz_5) begin
            tlbStorage_3_pp0_mat <= entryToFill_pp0_mat;
          end
          if(_zz_2) begin
            tlbStorage_0_pp0_d <= entryToFill_pp0_d;
          end
          if(_zz_3) begin
            tlbStorage_1_pp0_d <= entryToFill_pp0_d;
          end
          if(_zz_4) begin
            tlbStorage_2_pp0_d <= entryToFill_pp0_d;
          end
          if(_zz_5) begin
            tlbStorage_3_pp0_d <= entryToFill_pp0_d;
          end
          if(_zz_2) begin
            tlbStorage_0_pp0_v <= entryToFill_pp0_v;
          end
          if(_zz_3) begin
            tlbStorage_1_pp0_v <= entryToFill_pp0_v;
          end
          if(_zz_4) begin
            tlbStorage_2_pp0_v <= entryToFill_pp0_v;
          end
          if(_zz_5) begin
            tlbStorage_3_pp0_v <= entryToFill_pp0_v;
          end
          if(_zz_2) begin
            tlbStorage_0_pp1_ppn <= entryToFill_pp1_ppn;
          end
          if(_zz_3) begin
            tlbStorage_1_pp1_ppn <= entryToFill_pp1_ppn;
          end
          if(_zz_4) begin
            tlbStorage_2_pp1_ppn <= entryToFill_pp1_ppn;
          end
          if(_zz_5) begin
            tlbStorage_3_pp1_ppn <= entryToFill_pp1_ppn;
          end
          if(_zz_2) begin
            tlbStorage_0_pp1_plv <= entryToFill_pp1_plv;
          end
          if(_zz_3) begin
            tlbStorage_1_pp1_plv <= entryToFill_pp1_plv;
          end
          if(_zz_4) begin
            tlbStorage_2_pp1_plv <= entryToFill_pp1_plv;
          end
          if(_zz_5) begin
            tlbStorage_3_pp1_plv <= entryToFill_pp1_plv;
          end
          if(_zz_2) begin
            tlbStorage_0_pp1_mat <= entryToFill_pp1_mat;
          end
          if(_zz_3) begin
            tlbStorage_1_pp1_mat <= entryToFill_pp1_mat;
          end
          if(_zz_4) begin
            tlbStorage_2_pp1_mat <= entryToFill_pp1_mat;
          end
          if(_zz_5) begin
            tlbStorage_3_pp1_mat <= entryToFill_pp1_mat;
          end
          if(_zz_2) begin
            tlbStorage_0_pp1_d <= entryToFill_pp1_d;
          end
          if(_zz_3) begin
            tlbStorage_1_pp1_d <= entryToFill_pp1_d;
          end
          if(_zz_4) begin
            tlbStorage_2_pp1_d <= entryToFill_pp1_d;
          end
          if(_zz_5) begin
            tlbStorage_3_pp1_d <= entryToFill_pp1_d;
          end
          if(_zz_2) begin
            tlbStorage_0_pp1_v <= entryToFill_pp1_v;
          end
          if(_zz_3) begin
            tlbStorage_1_pp1_v <= entryToFill_pp1_v;
          end
          if(_zz_4) begin
            tlbStorage_2_pp1_v <= entryToFill_pp1_v;
          end
          if(_zz_5) begin
            tlbStorage_3_pp1_v <= entryToFill_pp1_v;
          end
        end
        TLBOp_fill : begin
          if(_zz_7) begin
            tlbStorage_0_vppn <= entryToFill_vppn;
          end
          if(_zz_8) begin
            tlbStorage_1_vppn <= entryToFill_vppn;
          end
          if(_zz_9) begin
            tlbStorage_2_vppn <= entryToFill_vppn;
          end
          if(_zz_10) begin
            tlbStorage_3_vppn <= entryToFill_vppn;
          end
          if(_zz_7) begin
            tlbStorage_0_ps <= entryToFill_ps;
          end
          if(_zz_8) begin
            tlbStorage_1_ps <= entryToFill_ps;
          end
          if(_zz_9) begin
            tlbStorage_2_ps <= entryToFill_ps;
          end
          if(_zz_10) begin
            tlbStorage_3_ps <= entryToFill_ps;
          end
          if(_zz_7) begin
            tlbStorage_0_g <= entryToFill_g;
          end
          if(_zz_8) begin
            tlbStorage_1_g <= entryToFill_g;
          end
          if(_zz_9) begin
            tlbStorage_2_g <= entryToFill_g;
          end
          if(_zz_10) begin
            tlbStorage_3_g <= entryToFill_g;
          end
          if(_zz_7) begin
            tlbStorage_0_asid <= entryToFill_asid;
          end
          if(_zz_8) begin
            tlbStorage_1_asid <= entryToFill_asid;
          end
          if(_zz_9) begin
            tlbStorage_2_asid <= entryToFill_asid;
          end
          if(_zz_10) begin
            tlbStorage_3_asid <= entryToFill_asid;
          end
          if(_zz_7) begin
            tlbStorage_0_e <= entryToFill_e;
          end
          if(_zz_8) begin
            tlbStorage_1_e <= entryToFill_e;
          end
          if(_zz_9) begin
            tlbStorage_2_e <= entryToFill_e;
          end
          if(_zz_10) begin
            tlbStorage_3_e <= entryToFill_e;
          end
          if(_zz_7) begin
            tlbStorage_0_pp0_ppn <= entryToFill_pp0_ppn;
          end
          if(_zz_8) begin
            tlbStorage_1_pp0_ppn <= entryToFill_pp0_ppn;
          end
          if(_zz_9) begin
            tlbStorage_2_pp0_ppn <= entryToFill_pp0_ppn;
          end
          if(_zz_10) begin
            tlbStorage_3_pp0_ppn <= entryToFill_pp0_ppn;
          end
          if(_zz_7) begin
            tlbStorage_0_pp0_plv <= entryToFill_pp0_plv;
          end
          if(_zz_8) begin
            tlbStorage_1_pp0_plv <= entryToFill_pp0_plv;
          end
          if(_zz_9) begin
            tlbStorage_2_pp0_plv <= entryToFill_pp0_plv;
          end
          if(_zz_10) begin
            tlbStorage_3_pp0_plv <= entryToFill_pp0_plv;
          end
          if(_zz_7) begin
            tlbStorage_0_pp0_mat <= entryToFill_pp0_mat;
          end
          if(_zz_8) begin
            tlbStorage_1_pp0_mat <= entryToFill_pp0_mat;
          end
          if(_zz_9) begin
            tlbStorage_2_pp0_mat <= entryToFill_pp0_mat;
          end
          if(_zz_10) begin
            tlbStorage_3_pp0_mat <= entryToFill_pp0_mat;
          end
          if(_zz_7) begin
            tlbStorage_0_pp0_d <= entryToFill_pp0_d;
          end
          if(_zz_8) begin
            tlbStorage_1_pp0_d <= entryToFill_pp0_d;
          end
          if(_zz_9) begin
            tlbStorage_2_pp0_d <= entryToFill_pp0_d;
          end
          if(_zz_10) begin
            tlbStorage_3_pp0_d <= entryToFill_pp0_d;
          end
          if(_zz_7) begin
            tlbStorage_0_pp0_v <= entryToFill_pp0_v;
          end
          if(_zz_8) begin
            tlbStorage_1_pp0_v <= entryToFill_pp0_v;
          end
          if(_zz_9) begin
            tlbStorage_2_pp0_v <= entryToFill_pp0_v;
          end
          if(_zz_10) begin
            tlbStorage_3_pp0_v <= entryToFill_pp0_v;
          end
          if(_zz_7) begin
            tlbStorage_0_pp1_ppn <= entryToFill_pp1_ppn;
          end
          if(_zz_8) begin
            tlbStorage_1_pp1_ppn <= entryToFill_pp1_ppn;
          end
          if(_zz_9) begin
            tlbStorage_2_pp1_ppn <= entryToFill_pp1_ppn;
          end
          if(_zz_10) begin
            tlbStorage_3_pp1_ppn <= entryToFill_pp1_ppn;
          end
          if(_zz_7) begin
            tlbStorage_0_pp1_plv <= entryToFill_pp1_plv;
          end
          if(_zz_8) begin
            tlbStorage_1_pp1_plv <= entryToFill_pp1_plv;
          end
          if(_zz_9) begin
            tlbStorage_2_pp1_plv <= entryToFill_pp1_plv;
          end
          if(_zz_10) begin
            tlbStorage_3_pp1_plv <= entryToFill_pp1_plv;
          end
          if(_zz_7) begin
            tlbStorage_0_pp1_mat <= entryToFill_pp1_mat;
          end
          if(_zz_8) begin
            tlbStorage_1_pp1_mat <= entryToFill_pp1_mat;
          end
          if(_zz_9) begin
            tlbStorage_2_pp1_mat <= entryToFill_pp1_mat;
          end
          if(_zz_10) begin
            tlbStorage_3_pp1_mat <= entryToFill_pp1_mat;
          end
          if(_zz_7) begin
            tlbStorage_0_pp1_d <= entryToFill_pp1_d;
          end
          if(_zz_8) begin
            tlbStorage_1_pp1_d <= entryToFill_pp1_d;
          end
          if(_zz_9) begin
            tlbStorage_2_pp1_d <= entryToFill_pp1_d;
          end
          if(_zz_10) begin
            tlbStorage_3_pp1_d <= entryToFill_pp1_d;
          end
          if(_zz_7) begin
            tlbStorage_0_pp1_v <= entryToFill_pp1_v;
          end
          if(_zz_8) begin
            tlbStorage_1_pp1_v <= entryToFill_pp1_v;
          end
          if(_zz_9) begin
            tlbStorage_2_pp1_v <= entryToFill_pp1_v;
          end
          if(_zz_10) begin
            tlbStorage_3_pp1_v <= entryToFill_pp1_v;
          end
        end
        TLBOp_inv : begin
          if(when_TLB_l130) begin
            if(_zz_11[0]) begin
              tlbStorage_0_e <= 1'b0;
            end
            if(_zz_11[1]) begin
              tlbStorage_1_e <= 1'b0;
            end
            if(_zz_11[2]) begin
              tlbStorage_2_e <= 1'b0;
            end
            if(_zz_11[3]) begin
              tlbStorage_3_e <= 1'b0;
            end
          end
        end
        default : begin
        end
      endcase
    end
  end


endmodule

module AXIArbiter (
  output wire [3:0]    io_out_arid,
  output wire [31:0]   io_out_araddr,
  output wire [7:0]    io_out_arlen,
  output wire [2:0]    io_out_arsize,
  output wire [1:0]    io_out_arburst,
  output wire [1:0]    io_out_arlock,
  output wire [3:0]    io_out_arcache,
  output wire [2:0]    io_out_arprot,
  output wire          io_out_arvalid,
  input  wire          io_out_arready,
  input  wire [3:0]    io_out_rid,
  input  wire [31:0]   io_out_rdata,
  input  wire [1:0]    io_out_rresp,
  input  wire          io_out_rlast,
  input  wire          io_out_rvalid,
  output wire          io_out_rready,
  output wire [3:0]    io_out_awid,
  output wire [31:0]   io_out_awaddr,
  output wire [7:0]    io_out_awlen,
  output wire [2:0]    io_out_awsize,
  output wire [1:0]    io_out_awburst,
  output wire [1:0]    io_out_awlock,
  output wire [3:0]    io_out_awcache,
  output wire [2:0]    io_out_awprot,
  output wire          io_out_awvalid,
  input  wire          io_out_awready,
  output wire [3:0]    io_out_wid,
  output wire [31:0]   io_out_wdata,
  output wire [3:0]    io_out_wstrb,
  output wire          io_out_wlast,
  output wire          io_out_wvalid,
  input  wire          io_out_wready,
  input  wire [3:0]    io_out_bid,
  input  wire [1:0]    io_out_bresp,
  input  wire          io_out_bvalid,
  output wire          io_out_bready,
  input  wire [3:0]    io_iCache_arid,
  input  wire [31:0]   io_iCache_araddr,
  input  wire [7:0]    io_iCache_arlen,
  input  wire [2:0]    io_iCache_arsize,
  input  wire [1:0]    io_iCache_arburst,
  input  wire [1:0]    io_iCache_arlock,
  input  wire [3:0]    io_iCache_arcache,
  input  wire [2:0]    io_iCache_arprot,
  input  wire          io_iCache_arvalid,
  output wire          io_iCache_arready,
  output wire [3:0]    io_iCache_rid,
  output wire [31:0]   io_iCache_rdata,
  output wire [1:0]    io_iCache_rresp,
  output wire          io_iCache_rlast,
  output wire          io_iCache_rvalid,
  input  wire          io_iCache_rready,
  input  wire [3:0]    io_dCache_arid,
  input  wire [31:0]   io_dCache_araddr,
  input  wire [7:0]    io_dCache_arlen,
  input  wire [2:0]    io_dCache_arsize,
  input  wire [1:0]    io_dCache_arburst,
  input  wire [1:0]    io_dCache_arlock,
  input  wire [3:0]    io_dCache_arcache,
  input  wire [2:0]    io_dCache_arprot,
  input  wire          io_dCache_arvalid,
  output wire          io_dCache_arready,
  output wire [3:0]    io_dCache_rid,
  output wire [31:0]   io_dCache_rdata,
  output wire [1:0]    io_dCache_rresp,
  output wire          io_dCache_rlast,
  output wire          io_dCache_rvalid,
  input  wire          io_dCache_rready,
  input  wire [3:0]    io_dCache_awid,
  input  wire [31:0]   io_dCache_awaddr,
  input  wire [7:0]    io_dCache_awlen,
  input  wire [2:0]    io_dCache_awsize,
  input  wire [1:0]    io_dCache_awburst,
  input  wire [1:0]    io_dCache_awlock,
  input  wire [3:0]    io_dCache_awcache,
  input  wire [2:0]    io_dCache_awprot,
  input  wire          io_dCache_awvalid,
  output wire          io_dCache_awready,
  input  wire [3:0]    io_dCache_wid,
  input  wire [31:0]   io_dCache_wdata,
  input  wire [3:0]    io_dCache_wstrb,
  input  wire          io_dCache_wlast,
  input  wire          io_dCache_wvalid,
  output wire          io_dCache_wready,
  output wire [3:0]    io_dCache_bid,
  output wire [1:0]    io_dCache_bresp,
  output wire          io_dCache_bvalid,
  input  wire          io_dCache_bready
);

  wire       [3:0]    _zz_chooseDCacheR;
  wire       [0:0]    _zz_chooseDCacheR_1;
  wire                chooseDCacheR;

  assign _zz_chooseDCacheR_1 = 1'b1;
  assign _zz_chooseDCacheR = {3'd0, _zz_chooseDCacheR_1};
  assign chooseDCacheR = (io_out_rid == _zz_chooseDCacheR);
  assign io_out_arid = (io_dCache_arvalid ? io_dCache_arid : io_iCache_arid);
  assign io_out_araddr = (io_dCache_arvalid ? io_dCache_araddr : io_iCache_araddr);
  assign io_out_arlen = (io_dCache_arvalid ? io_dCache_arlen : io_iCache_arlen);
  assign io_out_arsize = (io_dCache_arvalid ? io_dCache_arsize : io_iCache_arsize);
  assign io_out_arburst = (io_dCache_arvalid ? io_dCache_arburst : io_iCache_arburst);
  assign io_out_arlock = (io_dCache_arvalid ? io_dCache_arlock : io_iCache_arlock);
  assign io_out_arcache = (io_dCache_arvalid ? io_dCache_arcache : io_iCache_arcache);
  assign io_out_arprot = (io_dCache_arvalid ? io_dCache_arprot : io_iCache_arprot);
  assign io_out_arvalid = (io_dCache_arvalid ? io_dCache_arvalid : io_iCache_arvalid);
  assign io_iCache_arready = (io_out_arready && (! io_dCache_arvalid));
  assign io_dCache_arready = (io_out_arready && io_dCache_arvalid);
  assign io_iCache_rid = io_out_rid;
  assign io_iCache_rdata = io_out_rdata;
  assign io_iCache_rresp = io_out_rresp;
  assign io_iCache_rlast = io_out_rlast;
  assign io_iCache_rvalid = (io_out_rvalid && (! chooseDCacheR));
  assign io_dCache_rid = io_out_rid;
  assign io_dCache_rdata = io_out_rdata;
  assign io_dCache_rresp = io_out_rresp;
  assign io_dCache_rlast = io_out_rlast;
  assign io_dCache_rvalid = (io_out_rvalid && chooseDCacheR);
  assign io_out_rready = (chooseDCacheR ? io_dCache_rready : io_iCache_rready);
  assign io_out_awid = io_dCache_awid;
  assign io_out_awaddr = io_dCache_awaddr;
  assign io_out_awlen = io_dCache_awlen;
  assign io_out_awsize = io_dCache_awsize;
  assign io_out_awburst = io_dCache_awburst;
  assign io_out_awlock = io_dCache_awlock;
  assign io_out_awcache = io_dCache_awcache;
  assign io_out_awprot = io_dCache_awprot;
  assign io_out_awvalid = io_dCache_awvalid;
  assign io_dCache_awready = io_out_awready;
  assign io_out_wid = io_dCache_wid;
  assign io_out_wdata = io_dCache_wdata;
  assign io_out_wstrb = io_dCache_wstrb;
  assign io_out_wlast = io_dCache_wlast;
  assign io_out_wvalid = io_dCache_wvalid;
  assign io_dCache_wready = io_out_wready;
  assign io_dCache_bid = io_out_bid;
  assign io_dCache_bresp = io_out_bresp;
  assign io_dCache_bvalid = io_out_bready;
  assign io_out_bready = io_dCache_bready;

endmodule

//Decoder_1 replaced by Decoder

module Decoder (
  input  wire [31:0]   io_info_inst,
  input  wire [31:0]   io_info_branchInfo_predictPC,
  input  wire          io_info_branchInfo_predictResult,
  input  wire          io_info_exceptionInfo_exception,
  input  wire [5:0]    io_info_exceptionInfo_eCode,
  input  wire [0:0]    io_info_exceptionInfo_eSubCode,
  input  wire [31:0]   io_info_pc,
  input  wire [1:0]    _zz_when_Decoder_l40,
  output wire [31:0]   io_branchInfo_predictPC,
  output wire          io_branchInfo_predictResult,
  output wire [31:0]   io_branchResult_targetPC,
  output wire          io_branchResult_branchResult,
  output wire          io_branchResult_predictFail,
  output reg           io_exceptionInfo_exception,
  output reg  [5:0]    io_exceptionInfo_eCode,
  output reg  [0:0]    io_exceptionInfo_eSubCode,
  output wire [31:0]   io_pc,
  output reg  [3:0]    io_specialOp,
  output reg  [31:0]   io_imm,
  output reg  [3:0]    io_uopALU0_aluOp,
  output reg  [1:0]    io_uopALU0_bruOp,
  output reg  [1:0]    io_uopALU0_cruOp,
  output reg  [3:0]    io_uopALU1_aluOp,
  output reg  [1:0]    io_uopALU1_bruOp,
  output reg  [1:0]    io_uopMULU_muluOp,
  output reg  [1:0]    io_uopDIVU_divuOp,
  output reg  [3:0]    io_uopLSU_lsuOp,
  output reg  [4:0]    io_uopLSU_lsuCoOp,
  output reg  [2:0]    io_roopALU0_aluROOp,
  output reg  [2:0]    io_roopALU1_aluROOp,
  output reg  [1:0]    io_roopALU1_cruROOp,
  output reg  [0:0]    io_roopLSU_lsuROOp
);
  localparam ROBSpecialOp_nop = 4'd0;
  localparam ROBSpecialOp_bpuUpdate = 4'd1;
  localparam ROBSpecialOp_lsuAction = 4'd2;
  localparam ROBSpecialOp_ll = 4'd3;
  localparam ROBSpecialOp_writeCSR = 4'd4;
  localparam ROBSpecialOp_ertn = 4'd5;
  localparam ROBSpecialOp_idle = 4'd6;
  localparam ROBSpecialOp_readCSR = 4'd7;
  localparam ROBSpecialOp_readCNT = 4'd8;
  localparam ALUOp_add = 4'd0;
  localparam ALUOp_sub = 4'd1;
  localparam ALUOp_slt = 4'd2;
  localparam ALUOp_sltu = 4'd3;
  localparam ALUOp_eq = 4'd4;
  localparam ALUOp_nor_1 = 4'd5;
  localparam ALUOp_and_1 = 4'd6;
  localparam ALUOp_or_1 = 4'd7;
  localparam ALUOp_xor_1 = 4'd8;
  localparam ALUOp_sll_1 = 4'd9;
  localparam ALUOp_srl_1 = 4'd10;
  localparam ALUOp_sra_1 = 4'd11;
  localparam ALUOp_passa = 4'd12;
  localparam ALUOp_passb = 4'd13;
  localparam BRUOp_nop = 2'd0;
  localparam BRUOp_add = 2'd1;
  localparam BRUOp_cadd = 2'd2;
  localparam BRUOp_ncadd = 2'd3;
  localparam CRUOp_nop = 2'd0;
  localparam CRUOp_pass = 2'd1;
  localparam CRUOp_mask = 2'd2;
  localparam MULUOp_mullo = 2'd0;
  localparam MULUOp_mulhi = 2'd1;
  localparam MULUOp_mulhiu = 2'd2;
  localparam DIVUOp_div = 2'd0;
  localparam DIVUOp_divu = 2'd1;
  localparam DIVUOp_mod_1 = 2'd2;
  localparam DIVUOp_modu = 2'd3;
  localparam LSUOp_cacop = 4'd0;
  localparam LSUOp_tlbsrch = 4'd1;
  localparam LSUOp_tlbrd = 4'd2;
  localparam LSUOp_tlbwr = 4'd3;
  localparam LSUOp_tlbfill = 4'd4;
  localparam LSUOp_invtlb = 4'd5;
  localparam LSUOp_ll = 4'd6;
  localparam LSUOp_sc = 4'd7;
  localparam LSUOp_ld = 4'd8;
  localparam LSUOp_ldu = 4'd9;
  localparam LSUOp_st = 4'd10;
  localparam LSUOp_preld = 4'd11;
  localparam LSUOp_dbar = 4'd12;
  localparam LSUOp_ibar = 4'd13;
  localparam ALUROOp_reg_1 = 3'd0;
  localparam ALUROOp_regimm = 3'd1;
  localparam ALUROOp_pcimm = 3'd2;
  localparam ALUROOp_csr = 3'd3;
  localparam ALUROOp_linkpc = 3'd4;
  localparam ALUROOp_linkreg = 3'd5;
  localparam CRUROOp_id = 2'd0;
  localparam CRUROOp_lo = 2'd1;
  localparam CRUROOp_hi = 2'd2;
  localparam LSUROOp_reg_1 = 1'd0;
  localparam LSUROOp_regimm = 1'd1;
  localparam LSUSizeOp_byte_1 = 4'd1;
  localparam LSUSizeOp_halfword = 4'd3;
  localparam LSUSizeOp_word = 4'd15;

  wire       [3:0]    _zz_io_exceptionInfo_eCode;
  wire       [3:0]    _zz_io_exceptionInfo_eCode_1;
  wire       [3:0]    _zz_io_exceptionInfo_eCode_2;
  wire       [3:0]    _zz_io_exceptionInfo_eCode_3;
  wire       [0:0]    _zz_imm8_1;
  wire       [13:0]   _zz_imm8_2;
  wire       [0:0]    _zz_imm12_1;
  wire       [9:0]    _zz_imm12_2;
  wire       [0:0]    _zz_imm14_1;
  wire       [7:0]    _zz_imm14_2;
  wire       [0:0]    _zz_imm16_1;
  wire       [5:0]    _zz_imm16_2;
  wire       [0:0]    _zz_imm21_1;
  wire       [1:0]    _zz_imm21_2;
  wire       [31:0]   _zz_uimm5;
  wire       [4:0]    _zz_uimm5_1;
  wire       [31:0]   _zz_uimm12;
  wire       [11:0]   _zz_uimm12_1;
  wire       [31:0]   _zz_uimm14;
  wire       [13:0]   _zz_uimm14_1;
  wire       [4:0]    _zz_when_Decoder_l283;
  wire       [0:0]    _zz_when_Decoder_l283_1;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_10;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_11;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_12;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_13;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_14;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_15;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_16;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_17;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_18;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_19;
  reg                 privileged;
  reg                 illegal;
  reg                 break_1;
  reg                 syscall;
  wire                when_Decoder_l39;
  wire                when_Decoder_l40;
  wire                _zz_imm8;
  wire       [31:0]   imm8;
  wire                _zz_imm12;
  wire       [31:0]   imm12;
  wire                _zz_imm14;
  wire       [31:0]   imm14;
  wire                _zz_imm16;
  wire       [31:0]   imm16;
  wire                _zz_imm21;
  wire       [31:0]   imm21;
  wire                _zz_imm26;
  wire       [31:0]   imm26;
  wire       [31:0]   uimm5;
  wire       [31:0]   uimm12;
  wire       [31:0]   uimm14;
  wire       [31:0]   immu20;
  wire       [4:0]    lsuCoOp;
  wire                when_Decoder_l283;
  wire                when_Decoder_l285;
  wire                when_Decoder_l289;
  wire                when_Decoder_l294;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_1;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_2;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_3;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_4;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_5;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_6;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_7;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_8;
  wire       [3:0]    _zz_io_uopLSU_lsuCoOp_9;
  `ifndef SYNTHESIS
  reg [71:0] io_specialOp_string;
  reg [39:0] io_uopALU0_aluOp_string;
  reg [39:0] io_uopALU0_bruOp_string;
  reg [31:0] io_uopALU0_cruOp_string;
  reg [39:0] io_uopALU1_aluOp_string;
  reg [39:0] io_uopALU1_bruOp_string;
  reg [47:0] io_uopMULU_muluOp_string;
  reg [39:0] io_uopDIVU_divuOp_string;
  reg [55:0] io_uopLSU_lsuOp_string;
  reg [55:0] io_roopALU0_aluROOp_string;
  reg [55:0] io_roopALU1_aluROOp_string;
  reg [15:0] io_roopALU1_cruROOp_string;
  reg [47:0] io_roopLSU_lsuROOp_string;
  reg [63:0] _zz_io_uopLSU_lsuCoOp_string;
  reg [63:0] _zz_io_uopLSU_lsuCoOp_1_string;
  reg [63:0] _zz_io_uopLSU_lsuCoOp_2_string;
  reg [63:0] _zz_io_uopLSU_lsuCoOp_3_string;
  reg [63:0] _zz_io_uopLSU_lsuCoOp_4_string;
  reg [63:0] _zz_io_uopLSU_lsuCoOp_5_string;
  reg [63:0] _zz_io_uopLSU_lsuCoOp_6_string;
  reg [63:0] _zz_io_uopLSU_lsuCoOp_7_string;
  reg [63:0] _zz_io_uopLSU_lsuCoOp_8_string;
  reg [63:0] _zz_io_uopLSU_lsuCoOp_9_string;
  `endif


  assign _zz_io_exceptionInfo_eCode = 4'b1110;
  assign _zz_io_exceptionInfo_eCode_1 = 4'b1101;
  assign _zz_io_exceptionInfo_eCode_2 = 4'b1100;
  assign _zz_io_exceptionInfo_eCode_3 = 4'b1011;
  assign _zz_uimm5_1 = io_info_inst[14 : 10];
  assign _zz_uimm5 = {27'd0, _zz_uimm5_1};
  assign _zz_uimm12_1 = io_info_inst[21 : 10];
  assign _zz_uimm12 = {20'd0, _zz_uimm12_1};
  assign _zz_uimm14_1 = io_info_inst[23 : 10];
  assign _zz_uimm14 = {18'd0, _zz_uimm14_1};
  assign _zz_when_Decoder_l283_1 = 1'b1;
  assign _zz_when_Decoder_l283 = {4'd0, _zz_when_Decoder_l283_1};
  assign _zz_io_uopLSU_lsuCoOp_10 = _zz_io_uopLSU_lsuCoOp;
  assign _zz_io_uopLSU_lsuCoOp_11 = _zz_io_uopLSU_lsuCoOp_1;
  assign _zz_io_uopLSU_lsuCoOp_12 = _zz_io_uopLSU_lsuCoOp_2;
  assign _zz_io_uopLSU_lsuCoOp_13 = _zz_io_uopLSU_lsuCoOp_3;
  assign _zz_io_uopLSU_lsuCoOp_14 = _zz_io_uopLSU_lsuCoOp_4;
  assign _zz_io_uopLSU_lsuCoOp_15 = _zz_io_uopLSU_lsuCoOp_5;
  assign _zz_io_uopLSU_lsuCoOp_16 = _zz_io_uopLSU_lsuCoOp_6;
  assign _zz_io_uopLSU_lsuCoOp_17 = _zz_io_uopLSU_lsuCoOp_7;
  assign _zz_io_uopLSU_lsuCoOp_18 = _zz_io_uopLSU_lsuCoOp_8;
  assign _zz_io_uopLSU_lsuCoOp_19 = _zz_io_uopLSU_lsuCoOp_9;
  assign _zz_imm8_1 = _zz_imm8;
  assign _zz_imm8_2 = {_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,_zz_imm8}}}}}}}}}}}}};
  assign _zz_imm12_1 = _zz_imm12;
  assign _zz_imm12_2 = {_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,_zz_imm12}}}}}}}}};
  assign _zz_imm14_1 = _zz_imm14;
  assign _zz_imm14_2 = {_zz_imm14,{_zz_imm14,{_zz_imm14,{_zz_imm14,{_zz_imm14,{_zz_imm14,{_zz_imm14,_zz_imm14}}}}}}};
  assign _zz_imm16_1 = _zz_imm16;
  assign _zz_imm16_2 = {_zz_imm16,{_zz_imm16,{_zz_imm16,{_zz_imm16,{_zz_imm16,_zz_imm16}}}}};
  assign _zz_imm21_1 = _zz_imm21;
  assign _zz_imm21_2 = {_zz_imm21,_zz_imm21};
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_specialOp)
      ROBSpecialOp_nop : io_specialOp_string = "nop      ";
      ROBSpecialOp_bpuUpdate : io_specialOp_string = "bpuUpdate";
      ROBSpecialOp_lsuAction : io_specialOp_string = "lsuAction";
      ROBSpecialOp_ll : io_specialOp_string = "ll       ";
      ROBSpecialOp_writeCSR : io_specialOp_string = "writeCSR ";
      ROBSpecialOp_ertn : io_specialOp_string = "ertn     ";
      ROBSpecialOp_idle : io_specialOp_string = "idle     ";
      ROBSpecialOp_readCSR : io_specialOp_string = "readCSR  ";
      ROBSpecialOp_readCNT : io_specialOp_string = "readCNT  ";
      default : io_specialOp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_uopALU0_aluOp)
      ALUOp_add : io_uopALU0_aluOp_string = "add  ";
      ALUOp_sub : io_uopALU0_aluOp_string = "sub  ";
      ALUOp_slt : io_uopALU0_aluOp_string = "slt  ";
      ALUOp_sltu : io_uopALU0_aluOp_string = "sltu ";
      ALUOp_eq : io_uopALU0_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_uopALU0_aluOp_string = "nor_1";
      ALUOp_and_1 : io_uopALU0_aluOp_string = "and_1";
      ALUOp_or_1 : io_uopALU0_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_uopALU0_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_uopALU0_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_uopALU0_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_uopALU0_aluOp_string = "sra_1";
      ALUOp_passa : io_uopALU0_aluOp_string = "passa";
      ALUOp_passb : io_uopALU0_aluOp_string = "passb";
      default : io_uopALU0_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_uopALU0_bruOp)
      BRUOp_nop : io_uopALU0_bruOp_string = "nop  ";
      BRUOp_add : io_uopALU0_bruOp_string = "add  ";
      BRUOp_cadd : io_uopALU0_bruOp_string = "cadd ";
      BRUOp_ncadd : io_uopALU0_bruOp_string = "ncadd";
      default : io_uopALU0_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_uopALU0_cruOp)
      CRUOp_nop : io_uopALU0_cruOp_string = "nop ";
      CRUOp_pass : io_uopALU0_cruOp_string = "pass";
      CRUOp_mask : io_uopALU0_cruOp_string = "mask";
      default : io_uopALU0_cruOp_string = "????";
    endcase
  end
  always @(*) begin
    case(io_uopALU1_aluOp)
      ALUOp_add : io_uopALU1_aluOp_string = "add  ";
      ALUOp_sub : io_uopALU1_aluOp_string = "sub  ";
      ALUOp_slt : io_uopALU1_aluOp_string = "slt  ";
      ALUOp_sltu : io_uopALU1_aluOp_string = "sltu ";
      ALUOp_eq : io_uopALU1_aluOp_string = "eq   ";
      ALUOp_nor_1 : io_uopALU1_aluOp_string = "nor_1";
      ALUOp_and_1 : io_uopALU1_aluOp_string = "and_1";
      ALUOp_or_1 : io_uopALU1_aluOp_string = "or_1 ";
      ALUOp_xor_1 : io_uopALU1_aluOp_string = "xor_1";
      ALUOp_sll_1 : io_uopALU1_aluOp_string = "sll_1";
      ALUOp_srl_1 : io_uopALU1_aluOp_string = "srl_1";
      ALUOp_sra_1 : io_uopALU1_aluOp_string = "sra_1";
      ALUOp_passa : io_uopALU1_aluOp_string = "passa";
      ALUOp_passb : io_uopALU1_aluOp_string = "passb";
      default : io_uopALU1_aluOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_uopALU1_bruOp)
      BRUOp_nop : io_uopALU1_bruOp_string = "nop  ";
      BRUOp_add : io_uopALU1_bruOp_string = "add  ";
      BRUOp_cadd : io_uopALU1_bruOp_string = "cadd ";
      BRUOp_ncadd : io_uopALU1_bruOp_string = "ncadd";
      default : io_uopALU1_bruOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_uopMULU_muluOp)
      MULUOp_mullo : io_uopMULU_muluOp_string = "mullo ";
      MULUOp_mulhi : io_uopMULU_muluOp_string = "mulhi ";
      MULUOp_mulhiu : io_uopMULU_muluOp_string = "mulhiu";
      default : io_uopMULU_muluOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_uopDIVU_divuOp)
      DIVUOp_div : io_uopDIVU_divuOp_string = "div  ";
      DIVUOp_divu : io_uopDIVU_divuOp_string = "divu ";
      DIVUOp_mod_1 : io_uopDIVU_divuOp_string = "mod_1";
      DIVUOp_modu : io_uopDIVU_divuOp_string = "modu ";
      default : io_uopDIVU_divuOp_string = "?????";
    endcase
  end
  always @(*) begin
    case(io_uopLSU_lsuOp)
      LSUOp_cacop : io_uopLSU_lsuOp_string = "cacop  ";
      LSUOp_tlbsrch : io_uopLSU_lsuOp_string = "tlbsrch";
      LSUOp_tlbrd : io_uopLSU_lsuOp_string = "tlbrd  ";
      LSUOp_tlbwr : io_uopLSU_lsuOp_string = "tlbwr  ";
      LSUOp_tlbfill : io_uopLSU_lsuOp_string = "tlbfill";
      LSUOp_invtlb : io_uopLSU_lsuOp_string = "invtlb ";
      LSUOp_ll : io_uopLSU_lsuOp_string = "ll     ";
      LSUOp_sc : io_uopLSU_lsuOp_string = "sc     ";
      LSUOp_ld : io_uopLSU_lsuOp_string = "ld     ";
      LSUOp_ldu : io_uopLSU_lsuOp_string = "ldu    ";
      LSUOp_st : io_uopLSU_lsuOp_string = "st     ";
      LSUOp_preld : io_uopLSU_lsuOp_string = "preld  ";
      LSUOp_dbar : io_uopLSU_lsuOp_string = "dbar   ";
      LSUOp_ibar : io_uopLSU_lsuOp_string = "ibar   ";
      default : io_uopLSU_lsuOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_roopALU0_aluROOp)
      ALUROOp_reg_1 : io_roopALU0_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : io_roopALU0_aluROOp_string = "regimm ";
      ALUROOp_pcimm : io_roopALU0_aluROOp_string = "pcimm  ";
      ALUROOp_csr : io_roopALU0_aluROOp_string = "csr    ";
      ALUROOp_linkpc : io_roopALU0_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : io_roopALU0_aluROOp_string = "linkreg";
      default : io_roopALU0_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_roopALU1_aluROOp)
      ALUROOp_reg_1 : io_roopALU1_aluROOp_string = "reg_1  ";
      ALUROOp_regimm : io_roopALU1_aluROOp_string = "regimm ";
      ALUROOp_pcimm : io_roopALU1_aluROOp_string = "pcimm  ";
      ALUROOp_csr : io_roopALU1_aluROOp_string = "csr    ";
      ALUROOp_linkpc : io_roopALU1_aluROOp_string = "linkpc ";
      ALUROOp_linkreg : io_roopALU1_aluROOp_string = "linkreg";
      default : io_roopALU1_aluROOp_string = "???????";
    endcase
  end
  always @(*) begin
    case(io_roopALU1_cruROOp)
      CRUROOp_id : io_roopALU1_cruROOp_string = "id";
      CRUROOp_lo : io_roopALU1_cruROOp_string = "lo";
      CRUROOp_hi : io_roopALU1_cruROOp_string = "hi";
      default : io_roopALU1_cruROOp_string = "??";
    endcase
  end
  always @(*) begin
    case(io_roopLSU_lsuROOp)
      LSUROOp_reg_1 : io_roopLSU_lsuROOp_string = "reg_1 ";
      LSUROOp_regimm : io_roopLSU_lsuROOp_string = "regimm";
      default : io_roopLSU_lsuROOp_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_uopLSU_lsuCoOp)
      LSUSizeOp_byte_1 : _zz_io_uopLSU_lsuCoOp_string = "byte_1  ";
      LSUSizeOp_halfword : _zz_io_uopLSU_lsuCoOp_string = "halfword";
      LSUSizeOp_word : _zz_io_uopLSU_lsuCoOp_string = "word    ";
      default : _zz_io_uopLSU_lsuCoOp_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_uopLSU_lsuCoOp_1)
      LSUSizeOp_byte_1 : _zz_io_uopLSU_lsuCoOp_1_string = "byte_1  ";
      LSUSizeOp_halfword : _zz_io_uopLSU_lsuCoOp_1_string = "halfword";
      LSUSizeOp_word : _zz_io_uopLSU_lsuCoOp_1_string = "word    ";
      default : _zz_io_uopLSU_lsuCoOp_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_uopLSU_lsuCoOp_2)
      LSUSizeOp_byte_1 : _zz_io_uopLSU_lsuCoOp_2_string = "byte_1  ";
      LSUSizeOp_halfword : _zz_io_uopLSU_lsuCoOp_2_string = "halfword";
      LSUSizeOp_word : _zz_io_uopLSU_lsuCoOp_2_string = "word    ";
      default : _zz_io_uopLSU_lsuCoOp_2_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_uopLSU_lsuCoOp_3)
      LSUSizeOp_byte_1 : _zz_io_uopLSU_lsuCoOp_3_string = "byte_1  ";
      LSUSizeOp_halfword : _zz_io_uopLSU_lsuCoOp_3_string = "halfword";
      LSUSizeOp_word : _zz_io_uopLSU_lsuCoOp_3_string = "word    ";
      default : _zz_io_uopLSU_lsuCoOp_3_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_uopLSU_lsuCoOp_4)
      LSUSizeOp_byte_1 : _zz_io_uopLSU_lsuCoOp_4_string = "byte_1  ";
      LSUSizeOp_halfword : _zz_io_uopLSU_lsuCoOp_4_string = "halfword";
      LSUSizeOp_word : _zz_io_uopLSU_lsuCoOp_4_string = "word    ";
      default : _zz_io_uopLSU_lsuCoOp_4_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_uopLSU_lsuCoOp_5)
      LSUSizeOp_byte_1 : _zz_io_uopLSU_lsuCoOp_5_string = "byte_1  ";
      LSUSizeOp_halfword : _zz_io_uopLSU_lsuCoOp_5_string = "halfword";
      LSUSizeOp_word : _zz_io_uopLSU_lsuCoOp_5_string = "word    ";
      default : _zz_io_uopLSU_lsuCoOp_5_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_uopLSU_lsuCoOp_6)
      LSUSizeOp_byte_1 : _zz_io_uopLSU_lsuCoOp_6_string = "byte_1  ";
      LSUSizeOp_halfword : _zz_io_uopLSU_lsuCoOp_6_string = "halfword";
      LSUSizeOp_word : _zz_io_uopLSU_lsuCoOp_6_string = "word    ";
      default : _zz_io_uopLSU_lsuCoOp_6_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_uopLSU_lsuCoOp_7)
      LSUSizeOp_byte_1 : _zz_io_uopLSU_lsuCoOp_7_string = "byte_1  ";
      LSUSizeOp_halfword : _zz_io_uopLSU_lsuCoOp_7_string = "halfword";
      LSUSizeOp_word : _zz_io_uopLSU_lsuCoOp_7_string = "word    ";
      default : _zz_io_uopLSU_lsuCoOp_7_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_uopLSU_lsuCoOp_8)
      LSUSizeOp_byte_1 : _zz_io_uopLSU_lsuCoOp_8_string = "byte_1  ";
      LSUSizeOp_halfword : _zz_io_uopLSU_lsuCoOp_8_string = "halfword";
      LSUSizeOp_word : _zz_io_uopLSU_lsuCoOp_8_string = "word    ";
      default : _zz_io_uopLSU_lsuCoOp_8_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_uopLSU_lsuCoOp_9)
      LSUSizeOp_byte_1 : _zz_io_uopLSU_lsuCoOp_9_string = "byte_1  ";
      LSUSizeOp_halfword : _zz_io_uopLSU_lsuCoOp_9_string = "halfword";
      LSUSizeOp_word : _zz_io_uopLSU_lsuCoOp_9_string = "word    ";
      default : _zz_io_uopLSU_lsuCoOp_9_string = "????????";
    endcase
  end
  `endif

  always @(*) begin
    privileged = 1'b0;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
        privileged = 1'b1;
      end
      32'b0000011000?????????????????????? : begin
        if(when_Decoder_l294) begin
          privileged = 1'b1;
        end
      end
      32'b00000110010010000010100000000000 : begin
        privileged = 1'b1;
      end
      32'b00000110010010000010110000000000 : begin
        privileged = 1'b1;
      end
      32'b00000110010010000011000000000000 : begin
        privileged = 1'b1;
      end
      32'b00000110010010000011010000000000 : begin
        privileged = 1'b1;
      end
      32'b00000110010010000011100000000000 : begin
        privileged = 1'b1;
      end
      32'b00000110010010001??????????????? : begin
        privileged = 1'b1;
      end
      32'b00000110010010011??????????????? : begin
        privileged = 1'b1;
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110?????????????????????????? : begin
      end
      32'b010111?????????????????????????? : begin
      end
      32'b011000?????????????????????????? : begin
      end
      32'b011001?????????????????????????? : begin
      end
      32'b011010?????????????????????????? : begin
      end
      32'b011011?????????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    illegal = 1'b0;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110?????????????????????????? : begin
      end
      32'b010111?????????????????????????? : begin
      end
      32'b011000?????????????????????????? : begin
      end
      32'b011001?????????????????????????? : begin
      end
      32'b011010?????????????????????????? : begin
      end
      32'b011011?????????????????????????? : begin
      end
      default : begin
        illegal = 1'b1;
      end
    endcase
  end

  always @(*) begin
    break_1 = 1'b0;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
        break_1 = 1'b1;
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110?????????????????????????? : begin
      end
      32'b010111?????????????????????????? : begin
      end
      32'b011000?????????????????????????? : begin
      end
      32'b011001?????????????????????????? : begin
      end
      32'b011010?????????????????????????? : begin
      end
      32'b011011?????????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    syscall = 1'b0;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
        syscall = 1'b1;
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110?????????????????????????? : begin
      end
      32'b010111?????????????????????????? : begin
      end
      32'b011000?????????????????????????? : begin
      end
      32'b011001?????????????????????????? : begin
      end
      32'b011010?????????????????????????? : begin
      end
      32'b011011?????????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  assign when_Decoder_l39 = (! io_info_exceptionInfo_exception);
  assign when_Decoder_l40 = (privileged && (_zz_when_Decoder_l40 != 2'b00));
  always @(*) begin
    if(when_Decoder_l39) begin
      if(when_Decoder_l40) begin
        io_exceptionInfo_exception = 1'b1;
      end else begin
        if(illegal) begin
          io_exceptionInfo_exception = 1'b1;
        end else begin
          if(break_1) begin
            io_exceptionInfo_exception = 1'b1;
          end else begin
            if(syscall) begin
              io_exceptionInfo_exception = 1'b1;
            end else begin
              io_exceptionInfo_exception = io_info_exceptionInfo_exception;
            end
          end
        end
      end
    end else begin
      io_exceptionInfo_exception = io_info_exceptionInfo_exception;
    end
  end

  always @(*) begin
    if(when_Decoder_l39) begin
      if(when_Decoder_l40) begin
        io_exceptionInfo_eCode = {2'd0, _zz_io_exceptionInfo_eCode};
      end else begin
        if(illegal) begin
          io_exceptionInfo_eCode = {2'd0, _zz_io_exceptionInfo_eCode_1};
        end else begin
          if(break_1) begin
            io_exceptionInfo_eCode = {2'd0, _zz_io_exceptionInfo_eCode_2};
          end else begin
            if(syscall) begin
              io_exceptionInfo_eCode = {2'd0, _zz_io_exceptionInfo_eCode_3};
            end else begin
              io_exceptionInfo_eCode = io_info_exceptionInfo_eCode;
            end
          end
        end
      end
    end else begin
      io_exceptionInfo_eCode = io_info_exceptionInfo_eCode;
    end
  end

  always @(*) begin
    if(when_Decoder_l39) begin
      if(when_Decoder_l40) begin
        io_exceptionInfo_eSubCode = 1'b0;
      end else begin
        if(illegal) begin
          io_exceptionInfo_eSubCode = 1'b0;
        end else begin
          if(break_1) begin
            io_exceptionInfo_eSubCode = 1'b0;
          end else begin
            if(syscall) begin
              io_exceptionInfo_eSubCode = 1'b0;
            end else begin
              io_exceptionInfo_eSubCode = io_info_exceptionInfo_eSubCode;
            end
          end
        end
      end
    end else begin
      io_exceptionInfo_eSubCode = io_info_exceptionInfo_eSubCode;
    end
  end

  assign io_branchResult_targetPC = io_info_branchInfo_predictPC;
  assign io_branchResult_branchResult = 1'b0;
  assign io_branchResult_predictFail = io_info_branchInfo_predictResult;
  assign io_branchInfo_predictPC = io_info_branchInfo_predictPC;
  assign io_branchInfo_predictResult = io_info_branchInfo_predictResult;
  assign io_pc = io_info_pc;
  assign _zz_imm8 = io_info_inst[17];
  assign imm8 = {{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8,{_zz_imm8_1,_zz_imm8_2}}}}}}}}}},io_info_inst[17 : 10]};
  assign _zz_imm12 = io_info_inst[21];
  assign imm12 = {{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12,{_zz_imm12_1,_zz_imm12_2}}}}}}}}}},io_info_inst[21 : 10]};
  assign _zz_imm14 = io_info_inst[23];
  assign imm14 = ({{_zz_imm14,{_zz_imm14,{_zz_imm14,{_zz_imm14,{_zz_imm14,{_zz_imm14,{_zz_imm14,{_zz_imm14,{_zz_imm14,{_zz_imm14_1,_zz_imm14_2}}}}}}}}}},io_info_inst[23 : 10]} <<< 2);
  assign _zz_imm16 = io_info_inst[25];
  assign imm16 = {{_zz_imm16,{_zz_imm16,{_zz_imm16,{_zz_imm16,{_zz_imm16,{_zz_imm16,{_zz_imm16,{_zz_imm16,{_zz_imm16,{_zz_imm16_1,_zz_imm16_2}}}}}}}}}},io_info_inst[25 : 10]};
  assign _zz_imm21 = io_info_inst[4];
  assign imm21 = {{{_zz_imm21,{_zz_imm21,{_zz_imm21,{_zz_imm21,{_zz_imm21,{_zz_imm21,{_zz_imm21,{_zz_imm21,{_zz_imm21_1,_zz_imm21_2}}}}}}}}},io_info_inst[4 : 0]},io_info_inst[25 : 10]};
  assign _zz_imm26 = io_info_inst[9];
  assign imm26 = {{{_zz_imm26,{_zz_imm26,{_zz_imm26,{_zz_imm26,{_zz_imm26,_zz_imm26}}}}},io_info_inst[9 : 0]},io_info_inst[25 : 10]};
  assign uimm5 = _zz_uimm5;
  assign uimm12 = _zz_uimm12;
  assign uimm14 = _zz_uimm14;
  assign immu20 = {io_info_inst[24 : 5],12'h000};
  assign lsuCoOp = io_info_inst[4 : 0];
  always @(*) begin
    io_specialOp = ROBSpecialOp_nop;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
        io_specialOp = ROBSpecialOp_readCNT;
      end
      32'b000000000000000001100000000????? : begin
        io_specialOp = ROBSpecialOp_readCNT;
      end
      32'b000000000000000001100100000????? : begin
        io_specialOp = ROBSpecialOp_readCNT;
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
        if(when_Decoder_l289) begin
          io_specialOp = ROBSpecialOp_writeCSR;
        end
      end
      32'b0000011000?????????????????????? : begin
        io_specialOp = ROBSpecialOp_lsuAction;
      end
      32'b00000110010010000010100000000000 : begin
        io_specialOp = ROBSpecialOp_lsuAction;
      end
      32'b00000110010010000010110000000000 : begin
        io_specialOp = ROBSpecialOp_lsuAction;
      end
      32'b00000110010010000011000000000000 : begin
        io_specialOp = ROBSpecialOp_lsuAction;
      end
      32'b00000110010010000011010000000000 : begin
        io_specialOp = ROBSpecialOp_lsuAction;
      end
      32'b00000110010010000011100000000000 : begin
        io_specialOp = ROBSpecialOp_ertn;
      end
      32'b00000110010010001??????????????? : begin
        io_specialOp = ROBSpecialOp_idle;
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
        io_specialOp = ROBSpecialOp_ll;
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
        io_specialOp = ROBSpecialOp_lsuAction;
      end
      32'b010011?????????????????????????? : begin
        io_specialOp = ROBSpecialOp_bpuUpdate;
      end
      32'b010100?????????????????????????? : begin
        io_specialOp = ROBSpecialOp_bpuUpdate;
      end
      32'b010101?????????????????????????? : begin
        io_specialOp = ROBSpecialOp_bpuUpdate;
      end
      32'b010110?????????????????????????? : begin
        io_specialOp = ROBSpecialOp_bpuUpdate;
      end
      32'b010111?????????????????????????? : begin
        io_specialOp = ROBSpecialOp_bpuUpdate;
      end
      32'b011000?????????????????????????? : begin
        io_specialOp = ROBSpecialOp_bpuUpdate;
      end
      32'b011001?????????????????????????? : begin
        io_specialOp = ROBSpecialOp_bpuUpdate;
      end
      32'b011010?????????????????????????? : begin
        io_specialOp = ROBSpecialOp_bpuUpdate;
      end
      32'b011011?????????????????????????? : begin
        io_specialOp = ROBSpecialOp_bpuUpdate;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_imm = imm8;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
        io_imm = uimm5;
      end
      32'b00000000010001001??????????????? : begin
        io_imm = uimm5;
      end
      32'b00000000010010001??????????????? : begin
        io_imm = uimm5;
      end
      32'b0000001000?????????????????????? : begin
        io_imm = imm12;
      end
      32'b0000001001?????????????????????? : begin
        io_imm = imm12;
      end
      32'b0000001010?????????????????????? : begin
        io_imm = imm12;
      end
      32'b0000001101?????????????????????? : begin
        io_imm = uimm12;
      end
      32'b0000001110?????????????????????? : begin
        io_imm = uimm12;
      end
      32'b0000001111?????????????????????? : begin
        io_imm = uimm12;
      end
      32'b00000100???????????????????????? : begin
        io_imm = uimm14;
      end
      32'b0000011000?????????????????????? : begin
        io_imm = imm12;
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
        io_imm = immu20;
      end
      32'b0001110????????????????????????? : begin
        io_imm = immu20;
      end
      32'b00100000???????????????????????? : begin
        io_imm = imm14;
      end
      32'b00100001???????????????????????? : begin
        io_imm = imm14;
      end
      32'b0010100000?????????????????????? : begin
        io_imm = imm12;
      end
      32'b0010100001?????????????????????? : begin
        io_imm = imm12;
      end
      32'b0010100010?????????????????????? : begin
        io_imm = imm12;
      end
      32'b0010100100?????????????????????? : begin
        io_imm = imm12;
      end
      32'b0010100101?????????????????????? : begin
        io_imm = imm12;
      end
      32'b0010100110?????????????????????? : begin
        io_imm = imm12;
      end
      32'b0010101000?????????????????????? : begin
        io_imm = imm12;
      end
      32'b0010101001?????????????????????? : begin
        io_imm = imm12;
      end
      32'b0010101011?????????????????????? : begin
        io_imm = imm12;
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
        io_imm = imm16;
      end
      32'b010100?????????????????????????? : begin
        io_imm = imm26;
      end
      32'b010101?????????????????????????? : begin
        io_imm = imm26;
      end
      32'b010110?????????????????????????? : begin
        io_imm = imm16;
      end
      32'b010111?????????????????????????? : begin
        io_imm = imm16;
      end
      32'b011000?????????????????????????? : begin
        io_imm = imm16;
      end
      32'b011001?????????????????????????? : begin
        io_imm = imm16;
      end
      32'b011010?????????????????????????? : begin
        io_imm = imm16;
      end
      32'b011011?????????????????????????? : begin
        io_imm = imm16;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_uopALU0_aluOp = ALUOp_add;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
        io_uopALU0_aluOp = ALUOp_add;
      end
      32'b00000000000100010??????????????? : begin
        io_uopALU0_aluOp = ALUOp_sub;
      end
      32'b00000000000100100??????????????? : begin
        io_uopALU0_aluOp = ALUOp_slt;
      end
      32'b00000000000100101??????????????? : begin
        io_uopALU0_aluOp = ALUOp_sltu;
      end
      32'b00000000000101000??????????????? : begin
        io_uopALU0_aluOp = ALUOp_nor_1;
      end
      32'b00000000000101001??????????????? : begin
        io_uopALU0_aluOp = ALUOp_and_1;
      end
      32'b00000000000101010??????????????? : begin
        io_uopALU0_aluOp = ALUOp_or_1;
      end
      32'b00000000000101011??????????????? : begin
        io_uopALU0_aluOp = ALUOp_xor_1;
      end
      32'b00000000000101110??????????????? : begin
        io_uopALU0_aluOp = ALUOp_sll_1;
      end
      32'b00000000000101111??????????????? : begin
        io_uopALU0_aluOp = ALUOp_srl_1;
      end
      32'b00000000000110000??????????????? : begin
        io_uopALU0_aluOp = ALUOp_sra_1;
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
        io_uopALU0_aluOp = ALUOp_sll_1;
      end
      32'b00000000010001001??????????????? : begin
        io_uopALU0_aluOp = ALUOp_srl_1;
      end
      32'b00000000010010001??????????????? : begin
        io_uopALU0_aluOp = ALUOp_sra_1;
      end
      32'b0000001000?????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_slt;
      end
      32'b0000001001?????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_sltu;
      end
      32'b0000001010?????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_add;
      end
      32'b0000001101?????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_and_1;
      end
      32'b0000001110?????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_or_1;
      end
      32'b0000001111?????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_xor_1;
      end
      32'b00000100???????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_passa;
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_passb;
      end
      32'b0001110????????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_add;
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_add;
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_add;
      end
      32'b010110?????????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_eq;
      end
      32'b010111?????????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_eq;
      end
      32'b011000?????????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_slt;
      end
      32'b011001?????????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_slt;
      end
      32'b011010?????????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_sltu;
      end
      32'b011011?????????????????????????? : begin
        io_uopALU0_aluOp = ALUOp_sltu;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_uopALU0_bruOp = BRUOp_nop;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
        io_uopALU0_bruOp = BRUOp_add;
      end
      32'b010100?????????????????????????? : begin
        io_uopALU0_bruOp = BRUOp_add;
      end
      32'b010101?????????????????????????? : begin
        io_uopALU0_bruOp = BRUOp_add;
      end
      32'b010110?????????????????????????? : begin
        io_uopALU0_bruOp = BRUOp_cadd;
      end
      32'b010111?????????????????????????? : begin
        io_uopALU0_bruOp = BRUOp_ncadd;
      end
      32'b011000?????????????????????????? : begin
        io_uopALU0_bruOp = BRUOp_cadd;
      end
      32'b011001?????????????????????????? : begin
        io_uopALU0_bruOp = BRUOp_ncadd;
      end
      32'b011010?????????????????????????? : begin
        io_uopALU0_bruOp = BRUOp_cadd;
      end
      32'b011011?????????????????????????? : begin
        io_uopALU0_bruOp = BRUOp_ncadd;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_uopALU0_cruOp = CRUOp_nop;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
        if(when_Decoder_l283) begin
          io_uopALU0_cruOp = CRUOp_pass;
        end else begin
          if(when_Decoder_l285) begin
            io_uopALU0_cruOp = CRUOp_mask;
          end
        end
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110?????????????????????????? : begin
      end
      32'b010111?????????????????????????? : begin
      end
      32'b011000?????????????????????????? : begin
      end
      32'b011001?????????????????????????? : begin
      end
      32'b011010?????????????????????????? : begin
      end
      32'b011011?????????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_uopALU1_aluOp = ALUOp_add;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
        io_uopALU1_aluOp = ALUOp_passa;
      end
      32'b000000000000000001100000000????? : begin
        io_uopALU1_aluOp = ALUOp_passa;
      end
      32'b000000000000000001100100000????? : begin
        io_uopALU1_aluOp = ALUOp_passa;
      end
      32'b00000000000100000??????????????? : begin
        io_uopALU1_aluOp = ALUOp_add;
      end
      32'b00000000000100010??????????????? : begin
        io_uopALU1_aluOp = ALUOp_sub;
      end
      32'b00000000000100100??????????????? : begin
        io_uopALU1_aluOp = ALUOp_slt;
      end
      32'b00000000000100101??????????????? : begin
        io_uopALU1_aluOp = ALUOp_sltu;
      end
      32'b00000000000101000??????????????? : begin
        io_uopALU1_aluOp = ALUOp_nor_1;
      end
      32'b00000000000101001??????????????? : begin
        io_uopALU1_aluOp = ALUOp_and_1;
      end
      32'b00000000000101010??????????????? : begin
        io_uopALU1_aluOp = ALUOp_or_1;
      end
      32'b00000000000101011??????????????? : begin
        io_uopALU1_aluOp = ALUOp_xor_1;
      end
      32'b00000000000101110??????????????? : begin
        io_uopALU1_aluOp = ALUOp_sll_1;
      end
      32'b00000000000101111??????????????? : begin
        io_uopALU1_aluOp = ALUOp_srl_1;
      end
      32'b00000000000110000??????????????? : begin
        io_uopALU1_aluOp = ALUOp_sra_1;
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
        io_uopALU1_aluOp = ALUOp_sll_1;
      end
      32'b00000000010001001??????????????? : begin
        io_uopALU1_aluOp = ALUOp_srl_1;
      end
      32'b00000000010010001??????????????? : begin
        io_uopALU1_aluOp = ALUOp_sra_1;
      end
      32'b0000001000?????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_slt;
      end
      32'b0000001001?????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_sltu;
      end
      32'b0000001010?????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_add;
      end
      32'b0000001101?????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_and_1;
      end
      32'b0000001110?????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_or_1;
      end
      32'b0000001111?????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_xor_1;
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_passb;
      end
      32'b0001110????????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_add;
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_add;
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_add;
      end
      32'b010110?????????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_eq;
      end
      32'b010111?????????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_eq;
      end
      32'b011000?????????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_slt;
      end
      32'b011001?????????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_slt;
      end
      32'b011010?????????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_sltu;
      end
      32'b011011?????????????????????????? : begin
        io_uopALU1_aluOp = ALUOp_sltu;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_uopALU1_bruOp = BRUOp_nop;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
        io_uopALU1_bruOp = BRUOp_add;
      end
      32'b010100?????????????????????????? : begin
        io_uopALU1_bruOp = BRUOp_add;
      end
      32'b010101?????????????????????????? : begin
        io_uopALU1_bruOp = BRUOp_add;
      end
      32'b010110?????????????????????????? : begin
        io_uopALU1_bruOp = BRUOp_cadd;
      end
      32'b010111?????????????????????????? : begin
        io_uopALU1_bruOp = BRUOp_ncadd;
      end
      32'b011000?????????????????????????? : begin
        io_uopALU1_bruOp = BRUOp_cadd;
      end
      32'b011001?????????????????????????? : begin
        io_uopALU1_bruOp = BRUOp_ncadd;
      end
      32'b011010?????????????????????????? : begin
        io_uopALU1_bruOp = BRUOp_cadd;
      end
      32'b011011?????????????????????????? : begin
        io_uopALU1_bruOp = BRUOp_ncadd;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_uopMULU_muluOp = MULUOp_mullo;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
        io_uopMULU_muluOp = MULUOp_mullo;
      end
      32'b00000000000111001??????????????? : begin
        io_uopMULU_muluOp = MULUOp_mulhi;
      end
      32'b00000000000111010??????????????? : begin
        io_uopMULU_muluOp = MULUOp_mulhiu;
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110?????????????????????????? : begin
      end
      32'b010111?????????????????????????? : begin
      end
      32'b011000?????????????????????????? : begin
      end
      32'b011001?????????????????????????? : begin
      end
      32'b011010?????????????????????????? : begin
      end
      32'b011011?????????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_uopDIVU_divuOp = DIVUOp_div;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
        io_uopDIVU_divuOp = DIVUOp_div;
      end
      32'b00000000001000001??????????????? : begin
        io_uopDIVU_divuOp = DIVUOp_mod_1;
      end
      32'b00000000001000010??????????????? : begin
        io_uopDIVU_divuOp = DIVUOp_divu;
      end
      32'b00000000001000011??????????????? : begin
        io_uopDIVU_divuOp = DIVUOp_modu;
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110?????????????????????????? : begin
      end
      32'b010111?????????????????????????? : begin
      end
      32'b011000?????????????????????????? : begin
      end
      32'b011001?????????????????????????? : begin
      end
      32'b011010?????????????????????????? : begin
      end
      32'b011011?????????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_uopLSU_lsuOp = LSUOp_dbar;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_cacop;
      end
      32'b00000110010010000010100000000000 : begin
        io_uopLSU_lsuOp = LSUOp_tlbsrch;
      end
      32'b00000110010010000010110000000000 : begin
        io_uopLSU_lsuOp = LSUOp_tlbrd;
      end
      32'b00000110010010000011000000000000 : begin
        io_uopLSU_lsuOp = LSUOp_tlbwr;
      end
      32'b00000110010010000011010000000000 : begin
        io_uopLSU_lsuOp = LSUOp_tlbfill;
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
        io_uopLSU_lsuOp = LSUOp_invtlb;
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_ll;
      end
      32'b00100001???????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_sc;
      end
      32'b0010100000?????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_ld;
      end
      32'b0010100001?????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_ld;
      end
      32'b0010100010?????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_ld;
      end
      32'b0010100100?????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_st;
      end
      32'b0010100101?????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_st;
      end
      32'b0010100110?????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_st;
      end
      32'b0010101000?????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_ldu;
      end
      32'b0010101001?????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_ldu;
      end
      32'b0010101011?????????????????????? : begin
        io_uopLSU_lsuOp = LSUOp_preld;
      end
      32'b00111000011100100??????????????? : begin
        io_uopLSU_lsuOp = LSUOp_dbar;
      end
      32'b00111000011100101??????????????? : begin
        io_uopLSU_lsuOp = LSUOp_ibar;
      end
      32'b010011?????????????????????????? : begin
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110?????????????????????????? : begin
      end
      32'b010111?????????????????????????? : begin
      end
      32'b011000?????????????????????????? : begin
      end
      32'b011001?????????????????????????? : begin
      end
      32'b011010?????????????????????????? : begin
      end
      32'b011011?????????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_uopLSU_lsuCoOp = 5'h00;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
        io_uopLSU_lsuCoOp = lsuCoOp;
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
        io_uopLSU_lsuCoOp = lsuCoOp;
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
        io_uopLSU_lsuCoOp = {1'd0, _zz_io_uopLSU_lsuCoOp_10};
      end
      32'b00100001???????????????????????? : begin
        io_uopLSU_lsuCoOp = {1'd0, _zz_io_uopLSU_lsuCoOp_11};
      end
      32'b0010100000?????????????????????? : begin
        io_uopLSU_lsuCoOp = {1'd0, _zz_io_uopLSU_lsuCoOp_12};
      end
      32'b0010100001?????????????????????? : begin
        io_uopLSU_lsuCoOp = {1'd0, _zz_io_uopLSU_lsuCoOp_13};
      end
      32'b0010100010?????????????????????? : begin
        io_uopLSU_lsuCoOp = {1'd0, _zz_io_uopLSU_lsuCoOp_14};
      end
      32'b0010100100?????????????????????? : begin
        io_uopLSU_lsuCoOp = {1'd0, _zz_io_uopLSU_lsuCoOp_15};
      end
      32'b0010100101?????????????????????? : begin
        io_uopLSU_lsuCoOp = {1'd0, _zz_io_uopLSU_lsuCoOp_16};
      end
      32'b0010100110?????????????????????? : begin
        io_uopLSU_lsuCoOp = {1'd0, _zz_io_uopLSU_lsuCoOp_17};
      end
      32'b0010101000?????????????????????? : begin
        io_uopLSU_lsuCoOp = {1'd0, _zz_io_uopLSU_lsuCoOp_18};
      end
      32'b0010101001?????????????????????? : begin
        io_uopLSU_lsuCoOp = {1'd0, _zz_io_uopLSU_lsuCoOp_19};
      end
      32'b0010101011?????????????????????? : begin
        io_uopLSU_lsuCoOp = lsuCoOp;
      end
      32'b00111000011100100??????????????? : begin
        io_uopLSU_lsuCoOp = lsuCoOp;
      end
      32'b00111000011100101??????????????? : begin
        io_uopLSU_lsuCoOp = lsuCoOp;
      end
      32'b010011?????????????????????????? : begin
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110?????????????????????????? : begin
      end
      32'b010111?????????????????????????? : begin
      end
      32'b011000?????????????????????????? : begin
      end
      32'b011001?????????????????????????? : begin
      end
      32'b011010?????????????????????????? : begin
      end
      32'b011011?????????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_roopALU0_aluROOp = ALUROOp_reg_1;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000100010??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000100100??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000100101??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101000??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101001??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101010??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101011??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101110??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101111??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000110000??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_regimm;
      end
      32'b00000000010001001??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_regimm;
      end
      32'b00000000010010001??????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_regimm;
      end
      32'b0000001000?????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_regimm;
      end
      32'b0000001001?????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_regimm;
      end
      32'b0000001010?????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_regimm;
      end
      32'b0000001101?????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_regimm;
      end
      32'b0000001110?????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_regimm;
      end
      32'b0000001111?????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_regimm;
      end
      32'b00000100???????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_csr;
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_pcimm;
      end
      32'b0001110????????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_pcimm;
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_linkpc;
      end
      32'b010100?????????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b010101?????????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_linkreg;
      end
      32'b010110?????????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b010111?????????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b011000?????????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b011001?????????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b011010?????????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      32'b011011?????????????????????????? : begin
        io_roopALU0_aluROOp = ALUROOp_reg_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_roopALU1_aluROOp = ALUROOp_reg_1;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
        io_roopALU1_aluROOp = ALUROOp_csr;
      end
      32'b000000000000000001100000000????? : begin
        io_roopALU1_aluROOp = ALUROOp_csr;
      end
      32'b000000000000000001100100000????? : begin
        io_roopALU1_aluROOp = ALUROOp_csr;
      end
      32'b00000000000100000??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000100010??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000100100??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000100101??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101000??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101001??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101010??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101011??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101110??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000101111??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000110000??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_regimm;
      end
      32'b00000000010001001??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_regimm;
      end
      32'b00000000010010001??????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_regimm;
      end
      32'b0000001000?????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_regimm;
      end
      32'b0000001001?????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_regimm;
      end
      32'b0000001010?????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_regimm;
      end
      32'b0000001101?????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_regimm;
      end
      32'b0000001110?????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_regimm;
      end
      32'b0000001111?????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_regimm;
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_pcimm;
      end
      32'b0001110????????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_pcimm;
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_linkpc;
      end
      32'b010100?????????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b010101?????????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_linkreg;
      end
      32'b010110?????????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b010111?????????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b011000?????????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b011001?????????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b011010?????????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      32'b011011?????????????????????????? : begin
        io_roopALU1_aluROOp = ALUROOp_reg_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_roopALU1_cruROOp = CRUROOp_id;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
        io_roopALU1_cruROOp = CRUROOp_id;
      end
      32'b000000000000000001100000000????? : begin
        io_roopALU1_cruROOp = CRUROOp_lo;
      end
      32'b000000000000000001100100000????? : begin
        io_roopALU1_cruROOp = CRUROOp_hi;
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
      end
      32'b00000110010010000010100000000000 : begin
      end
      32'b00000110010010000010110000000000 : begin
      end
      32'b00000110010010000011000000000000 : begin
      end
      32'b00000110010010000011010000000000 : begin
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
      end
      32'b00100001???????????????????????? : begin
      end
      32'b0010100000?????????????????????? : begin
      end
      32'b0010100001?????????????????????? : begin
      end
      32'b0010100010?????????????????????? : begin
      end
      32'b0010100100?????????????????????? : begin
      end
      32'b0010100101?????????????????????? : begin
      end
      32'b0010100110?????????????????????? : begin
      end
      32'b0010101000?????????????????????? : begin
      end
      32'b0010101001?????????????????????? : begin
      end
      32'b0010101011?????????????????????? : begin
      end
      32'b00111000011100100??????????????? : begin
      end
      32'b00111000011100101??????????????? : begin
      end
      32'b010011?????????????????????????? : begin
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110?????????????????????????? : begin
      end
      32'b010111?????????????????????????? : begin
      end
      32'b011000?????????????????????????? : begin
      end
      32'b011001?????????????????????????? : begin
      end
      32'b011010?????????????????????????? : begin
      end
      32'b011011?????????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_roopLSU_lsuROOp = LSUROOp_regimm;
    casez(io_info_inst)
      32'b0000000000000000011000?????00000 : begin
      end
      32'b000000000000000001100000000????? : begin
      end
      32'b000000000000000001100100000????? : begin
      end
      32'b00000000000100000??????????????? : begin
      end
      32'b00000000000100010??????????????? : begin
      end
      32'b00000000000100100??????????????? : begin
      end
      32'b00000000000100101??????????????? : begin
      end
      32'b00000000000101000??????????????? : begin
      end
      32'b00000000000101001??????????????? : begin
      end
      32'b00000000000101010??????????????? : begin
      end
      32'b00000000000101011??????????????? : begin
      end
      32'b00000000000101110??????????????? : begin
      end
      32'b00000000000101111??????????????? : begin
      end
      32'b00000000000110000??????????????? : begin
      end
      32'b00000000000111000??????????????? : begin
      end
      32'b00000000000111001??????????????? : begin
      end
      32'b00000000000111010??????????????? : begin
      end
      32'b00000000001000000??????????????? : begin
      end
      32'b00000000001000001??????????????? : begin
      end
      32'b00000000001000010??????????????? : begin
      end
      32'b00000000001000011??????????????? : begin
      end
      32'b00000000001010100??????????????? : begin
      end
      32'b00000000001010110??????????????? : begin
      end
      32'b00000000010000001??????????????? : begin
      end
      32'b00000000010001001??????????????? : begin
      end
      32'b00000000010010001??????????????? : begin
      end
      32'b0000001000?????????????????????? : begin
      end
      32'b0000001001?????????????????????? : begin
      end
      32'b0000001010?????????????????????? : begin
      end
      32'b0000001101?????????????????????? : begin
      end
      32'b0000001110?????????????????????? : begin
      end
      32'b0000001111?????????????????????? : begin
      end
      32'b00000100???????????????????????? : begin
      end
      32'b0000011000?????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b00000110010010000010100000000000 : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b00000110010010000010110000000000 : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b00000110010010000011000000000000 : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b00000110010010000011010000000000 : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b00000110010010000011100000000000 : begin
      end
      32'b00000110010010001??????????????? : begin
      end
      32'b00000110010010011??????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_reg_1;
      end
      32'b0001010????????????????????????? : begin
      end
      32'b0001110????????????????????????? : begin
      end
      32'b00100000???????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b00100001???????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b0010100000?????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b0010100001?????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b0010100010?????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b0010100100?????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b0010100101?????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b0010100110?????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b0010101000?????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b0010101001?????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b0010101011?????????????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b00111000011100100??????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b00111000011100101??????????????? : begin
        io_roopLSU_lsuROOp = LSUROOp_regimm;
      end
      32'b010011?????????????????????????? : begin
      end
      32'b010100?????????????????????????? : begin
      end
      32'b010101?????????????????????????? : begin
      end
      32'b010110?????????????????????????? : begin
      end
      32'b010111?????????????????????????? : begin
      end
      32'b011000?????????????????????????? : begin
      end
      32'b011001?????????????????????????? : begin
      end
      32'b011010?????????????????????????? : begin
      end
      32'b011011?????????????????????????? : begin
      end
      default : begin
      end
    endcase
  end

  assign when_Decoder_l283 = (io_info_inst[9 : 5] == _zz_when_Decoder_l283);
  assign when_Decoder_l285 = (io_info_inst[9 : 5] != 5'h00);
  assign when_Decoder_l289 = (io_info_inst[9 : 5] != 5'h00);
  assign when_Decoder_l294 = (lsuCoOp[4 : 3] != 2'b10);
  assign _zz_io_uopLSU_lsuCoOp = LSUSizeOp_word;
  assign _zz_io_uopLSU_lsuCoOp_1 = LSUSizeOp_word;
  assign _zz_io_uopLSU_lsuCoOp_2 = LSUSizeOp_byte_1;
  assign _zz_io_uopLSU_lsuCoOp_3 = LSUSizeOp_halfword;
  assign _zz_io_uopLSU_lsuCoOp_4 = LSUSizeOp_word;
  assign _zz_io_uopLSU_lsuCoOp_5 = LSUSizeOp_byte_1;
  assign _zz_io_uopLSU_lsuCoOp_6 = LSUSizeOp_halfword;
  assign _zz_io_uopLSU_lsuCoOp_7 = LSUSizeOp_word;
  assign _zz_io_uopLSU_lsuCoOp_8 = LSUSizeOp_byte_1;
  assign _zz_io_uopLSU_lsuCoOp_9 = LSUSizeOp_halfword;

endmodule
